----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:12:54 05/19/2012 
-- Design Name: 
-- Module Name:    DSPtester - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_unsigned.all;
use IEEE.STD_LOGIC_ARITH.ALL;

Library UNISIM;
use UNISIM.vcomponents.all;

Library UNIMACRO;
use UNIMACRO.vcomponents.all; 


entity divisor is
    Port ( DATA_0_i : in  STD_LOGIC_VECTOR (11 downto 0);
           DATA_1_i : in  STD_LOGIC_VECTOR (11 downto 0);
           clk : in  STD_LOGIC;
           RESULT : out  STD_LOGIC_VECTOR (9 downto 0));
end divisor;

architecture Behavioral of divisor is

signal DATA_0 :  STD_LOGIC_VECTOR (11 downto 0);
signal DATA_1 :  STD_LOGIC_VECTOR (11 downto 0);

signal memDO : STD_LOGIC_VECTOR(35 DOWNTO 0):=X"FFFFFFFFF";
signal adr : STD_LOGIC_VECTOR(9 DOWNTO 0):="0000000001";
signal test2 : STD_LOGIC_VECTOR(35 DOWNTO 0);
signal test3 : STD_LOGIC_VECTOR(3 DOWNTO 0);

signal n1_sh : Integer range 0 to 16 :=0;
signal n0_sh : Integer range 0 to 16 :=0;
signal n01_sh : Integer range -64 to 64 :=10;
signal n01_sh_del : Integer range -64 to 64 :=10;

signal n_sh : Integer range -32 to 32 :=20;
signal shift_end : Integer range -64 to 64 :=20;
signal shift_end_del : Integer range -64 to 64 :=20;

signal DATA_0_n : STD_LOGIC_VECTOR(12 DOWNTO 0);
signal DATA_1_h_rs : STD_LOGIC_VECTOR(15 DOWNTO 0);
signal DATA_1_hml : STD_LOGIC_VECTOR(12 DOWNTO 0);
signal mult1 : STD_LOGIC_VECTOR(25 DOWNTO 0);
signal mult1_sh: STD_LOGIC_VECTOR(14 DOWNTO 0);
signal solution_us : STD_LOGIC_VECTOR(30 DOWNTO 0);
signal solution_us_del : STD_LOGIC_VECTOR(30 DOWNTO 0):= (others => '0');


begin

process (clk)

variable test : STD_LOGIC_VECTOR(39 DOWNTO 0) :=(others => '0');
variable DATA_1_h : STD_LOGIC_VECTOR(12 DOWNTO 0) :=(others => '0');
variable DATA_1_l : STD_LOGIC_VECTOR(12 DOWNTO 0) :=(others => '0');
variable DATA_1_n : STD_LOGIC_VECTOR(11 DOWNTO 0) :="101000101000";

begin
      if (clk'event and clk = '1') then


			DATA_0 <= DATA_0_i;					
			DATA_1 <= DATA_1_i + DATA_0_i;	


			--normalize Data_1 and save amount of shift steps necesarry
			if DATA_0  = "000000000000" then
				n1_sh <= 0;
				DATA_1_n := "000000000000";
			elsif (DATA_1(11) = '1') then
				n1_sh <= 0;
				DATA_1_n := DATA_1;
			elsif (DATA_1(10) = '1') then
				n1_sh <= 1;
				DATA_1_n := DATA_1(10 downto 0) & "0";
			elsif (DATA_1(9) = '1') then
				n1_sh <= 2;
				DATA_1_n := DATA_1(9 downto 0) & "00";
			elsif (DATA_1(8) = '1') then
				n1_sh <= 3;
				DATA_1_n := DATA_1(8 downto 0) & "000";
			elsif (DATA_1(7) = '1') then
				n1_sh <= 4;
				DATA_1_n := DATA_1(7 downto 0) & "0000";
			elsif (DATA_1(6) = '1') then
				n1_sh <= 5;
				DATA_1_n := DATA_1(6 downto 0) & "00000";
			elsif(DATA_1(5) = '1') then
				n1_sh <= 6;
				DATA_1_n := DATA_1(5 downto 0) & "000000";
			elsif (DATA_1(4) = '1') then
				n1_sh <= 7;
				DATA_1_n := DATA_1(4 downto 0) & "0000000";
			elsif(DATA_1(3) = '1') then
				n1_sh <= 8;
				DATA_1_n := DATA_1(3 downto 0) & "00000000";
			elsif(DATA_1(2) = '1') then
				n1_sh <= 9;
				DATA_1_n := DATA_1(2 downto 0) & "000000000";
			elsif(DATA_1(1) = '1') then
				n1_sh <= 10;
				DATA_1_n := DATA_1(1 downto 0) & "0000000000";
			elsif(DATA_1(0) = '1') then
				n1_sh <= 11;
				DATA_1_n := DATA_1(0) & "00000000000";
			end if;

			--normalize Data_0 and save amount of shift steps necesarry
			if DATA_0  = "000000000000" then
				n0_sh <= 0;
				DATA_0_n <= "0" & DATA_0;
			elsif (DATA_0(11) = '1') then
				n0_sh <= 0;
				DATA_0_n <= "0" & DATA_0;
			elsif (DATA_0(10) = '1') then
				n0_sh <= 1;
				DATA_0_n <= "0" & DATA_0(10 downto 0) & "0";
			elsif (DATA_0(9) = '1') then
				n0_sh <= 2;
				DATA_0_n <= "0" & DATA_0(9 downto 0) & "00";
			elsif (DATA_0(8) = '1') then
				n0_sh <= 3;
				DATA_0_n <= "0" & DATA_0(8 downto 0) & "000";
			elsif (DATA_0(7) = '1') then
				n0_sh <= 4;
				DATA_0_n <= "0" & DATA_0(7 downto 0) & "0000";
			elsif (DATA_0(6) = '1') then
				n0_sh <= 5;
				DATA_0_n <= "0" & DATA_0(6 downto 0) & "00000";
			elsif(DATA_0(5) = '1') then
				n0_sh <= 6;
				DATA_0_n <= "0" & DATA_0(5 downto 0) & "000000";
			elsif (DATA_0(4) = '1') then
				n0_sh <= 7;
				DATA_0_n <= "0" & DATA_0(4 downto 0) & "0000000";
			elsif(DATA_0(3) = '1') then
				n0_sh <= 8;
				DATA_0_n <= "0" & DATA_0(3 downto 0) & "00000000";
			elsif(DATA_0(2) = '1') then
				n0_sh <= 9;
				DATA_0_n <= "0" & DATA_0(2 downto 0) & "000000000";
			elsif(DATA_0(1) = '1') then
				n0_sh <= 10;
				DATA_0_n <= "0" & DATA_0(1 downto 0) & "0000000000";
			elsif(DATA_0(0) = '1') then
				n0_sh <= 11;
				DATA_0_n <= "0" & DATA_0(0) & "00000000000";
			end if;
			DATA_1_h := "0" & DATA_1_n(11 downto 6) & "000000"; --save upper 6 bits +sign bit in 13 bit vector
			DATA_1_l := "0000000" & DATA_1_n(5 downto 0);		 --save lower 6 bit  +sign bit in 13 bit vector
			adr <="0000" & DATA_1_n(11 downto 6);					 --set adresse for the lookup table
			DATA_1_hml <= DATA_1_h - DATA_1_l;						 --get difference of upper and lower bits, DATA_1_hml gets multiplied by DATA_0_n 


			n01_sh <= n0_sh-n1_sh;										 --get difference of shift steps necesarry to normalize denominator and divisor, n0 and n1 max shoulde be 11 => max=11, min=-11
			-- memDO <= BRAM(adr)
			-- multi1 <= DSP(DATA_1_hml * DATA_0_n)


			n01_sh_del <= n01_sh;										 --delay difference of shifts
			mult1_sh <= mult1(25 downto 11); 						 --save 14 bit result of DATA_1_hml * DATA_0_n (not 12 + 1SignBit because of possible error correction), gets multiplied by DATA_1_h_rs 
			DATA_1_h_rs<= "01" & memDO(13 downto 0);            --receive normalized reciproc square of DATA_1 from lookup, 0 is sign, 1 is not saved - normalization
			n_sh <= conv_integer(memDO(18 downto 14));          --receive shift steps of normalized reciproc square from lookup, max should be 24, min = 12


			shift_end <=n01_sh_del+ n_sh+1;                     --add all shift steps, max shoulde be 36 min=1
			-- solution_us <= DSP(mult1_sh * DATA_1_h_rs)

			
			solution_us_del <=solution_us;                      --delay, due to timing constraints in full design
			shift_end_del <= shift_end;								 --delay, due to timing constraints in full design


			test:="000000000" & solution_us_del;					 --9 zeros +1 sign zero, precision 10 bit
			if shift_end_del/=1 then
			Result <= test(shift_end_del-1 downto shift_end_del-10);--use shifts to get result
			else
			Result <="0000000000";
			end if;
		
		end if;

end process;

   MULT_MACRO_inst : MULT_MACRO
   generic map (
      DEVICE => "VIRTEX5",    -- Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6" 
      LATENCY => 1,           -- Desired clock cycle latency, 0-4
		WIDTH_A => 13,          -- Multiplier A-input bus width, 1-25 
      WIDTH_B => 13)          -- Multiplier B-input bus width, 1-18
   port map (
      P => mult1,     -- Multiplier ouput bus, width determined by WIDTH_P generic 
      A => DATA_1_hml,     -- Multiplier input A bus, width determined by WIDTH_A generic 
      B => Data_0_n,     -- Multiplier input B bus, width determined by WIDTH_B generic 
      CE => '1',   -- 1-bit active high input clock enable
      CLK => clk, -- 1-bit positive edge clock input
      RST => '0'  -- 1-bit input active high reset
   );

   MULT_MACRO_inst_1 : MULT_MACRO
   generic map (
      DEVICE => "VIRTEX5",    -- Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6" 
      LATENCY => 1,           -- Desired clock cycle latency, 0-4
		WIDTH_A =>15,          -- Multiplier A-input bus width, 1-25 
      WIDTH_B => 16)          -- Multiplier B-input bus width, 1-18
   port map (
      P => solution_us,     -- Multiplier ouput bus, width determined by WIDTH_P generic 
      A => mult1_sh,     -- Multiplier input A bus, width determined by WIDTH_A generic 
      B => DATA_1_h_rs,     -- Multiplier input B bus, width determined by WIDTH_B generic 
      CE => '1',   -- 1-bit active high input clock enable
      CLK => clk, -- 1-bit positive edge clock input
      RST => '0'  -- 1-bit input active high reset
   );


BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
 generic map (
    BRAM_SIZE => "36Kb", -- Target BRAM, "18Kb" or "36Kb" 
    DEVICE => "VIRTEX5", -- Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6" 
    DO_REG => 0, -- Optional output register (0 or 1)
    INIT => X"ABCDEFF12",   --  Initial values on output port
    INIT_FILE => "NONE",
    WRITE_WIDTH => 36,   -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
    READ_WIDTH => 36,   -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
    SIM_MODE => "FAST", -- Simulation: "SAFE" vs "FAST",                                        -- era SAFE
                        -- see "Synthesis and Simulation Design Guide" for details
    SRVAL => X"000000000",   -- Set/Reset value for port output
    WRITE_MODE => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE" 
    -- The following INIT_xx declarations specify the initial contents of the RAM

  	 INIT_00 => b"0000000000000101000100111001011100000000000001010011000111000111000000000000010011010001111010110000000000000100100000000000000000000000000001001011000111000111000000000000010000000000000000000000000000000011100000000000000000000000000000000000000000000000",
	 INIT_01 => b"0000000000000101100010001101000100000000000001011001001110010111000000000000010110100000111100100000000000000101101100011100011100000000000001010100001110110011000000000000010101010001111010110000000000000101011001010010001000000000000001010000000000000000",
	 INIT_02 => b"0000000000000110001110111110001000000000000001011100001110110011000000000000010111001010010011010000000000000101110100011110101100000000000001011101101011000101000000000000010111100101001000100000000000000101111100010110001000000000000001011000000000000000",
	 INIT_03 => b"0000000000000110000001000011001000000000000001100000100011010001000000000000011000001101111011010000000000000110000100111001011100000000000001100001100111100110000000000000011000100000111100100000000000000110001010001101101100000000000001100011000111000111",
	 INIT_04 => b"0000000000000110010101100010110000000000000001100101101011000101000000000000011001011111101111100000000000000110011001010010001000000000000001100110101011111111000000000000011001110001011000100000000000000110011110000101110000000000000001100000000000000000",
	 INIT_05 => b"0000000000000110101101101010101100000000000001101011101111100010000000000000011001000000101110100000000000000110010000111011001100000000000001100100011011100011000000000000011001001010010011010000000000000110010011011111100000000000000001100101000111101011",
	 INIT_06 => b"0000000000000110100101101010100000000000000001101001100111100110000000000000011010011101010100100000000000000110101000001111001000000000000001101010010011001001000000000000011010101000110110110000000000000110101011010010111000000000000001101011000111000111",
	 INIT_07 => b"0000000000000110100000100000110000000000000001101000010000110010000000000000011010000110011100110000000000000110100010001101000100000000000001101000101101001110000000000000011010001101111011010000000000000110100100001010111100000000000001101001001110010111",

	 INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

    INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
 
    INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",  

    INITP_08 => X"00000000000000000000000000000000000000000000000000000000000000FF",
    INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
    INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")


  port map (
    DO => memDO,      -- Output data
    ADDR => adr,  -- Input address
    CLK => 	clk,    -- Input clock
    DI => 	test2,      -- Input data port  
    EN =>	'1',      -- Input RAM enable
    REGCE => '0', -- Input output register enable
    RST => '0',    -- Input reset
    WE => test3       -- Input write enable
 );

			
end Behavioral;