----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:12:54 05/19/2012 
-- Design Name: 
-- Module Name:    DSPtester - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_unsigned.all;
use IEEE.STD_LOGIC_ARITH.ALL;

Library UNISIM;
use UNISIM.vcomponents.all;

Library UNIMACRO;
use UNIMACRO.vcomponents.all; 


entity divisor_15 is
    Port ( DATA_0_i : in  STD_LOGIC_VECTOR (14 downto 0);
           DATA_1_i : in  STD_LOGIC_VECTOR (14 downto 0);
           clk : in  STD_LOGIC;
           RESULT : out  STD_LOGIC_VECTOR (9 downto 0));
end divisor_15;

architecture Behavioral of divisor_15 is

signal DATA_0 :  STD_LOGIC_VECTOR (14 downto 0);
signal DATA_1 :  STD_LOGIC_VECTOR (14 downto 0);

signal memDO : STD_LOGIC_VECTOR(35 DOWNTO 0):=X"FFFFFFFFF";
signal memDO_B : STD_LOGIC_VECTOR(35 DOWNTO 0):=X"FFFFFFFFF";
signal adr : STD_LOGIC_VECTOR(9 DOWNTO 0):="0000000001";
signal adrB : STD_LOGIC_VECTOR(9 DOWNTO 0):="0000000001";
signal test2 : STD_LOGIC_VECTOR(35 DOWNTO 0);
signal test3 : STD_LOGIC_VECTOR(3 DOWNTO 0);

signal n1_sh : Integer range 0 to 16 :=0;
signal n0_sh : Integer range 0 to 16 :=0;
signal n01_sh : Integer range -64 to 64 :=10;
signal n01_sh_del : Integer range -64 to 64 :=10;

signal n_sh : Integer range 0 to 40 :=20;
signal shift_end : Integer range -64 to 64 :=20;
signal shift_end_del : Integer range -64 to 64 :=20;

signal DATA_0_n : STD_LOGIC_VECTOR(15 DOWNTO 0);
signal DATA_1_h_rs : STD_LOGIC_VECTOR(17 DOWNTO 0);
signal DATA_1_hml : STD_LOGIC_VECTOR(15 DOWNTO 0);
signal mult1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
signal mult1_sh: STD_LOGIC_VECTOR(16 DOWNTO 0);
signal solution_us : STD_LOGIC_VECTOR(34 DOWNTO 0);
signal solution_us_del : STD_LOGIC_VECTOR(34 DOWNTO 0):= (others => '0');


begin

process (clk)

variable test : STD_LOGIC_VECTOR(43 DOWNTO 0) :=(others => '0');
variable DATA_1_h : STD_LOGIC_VECTOR(15 DOWNTO 0) :=(others => '0');
variable DATA_1_l : STD_LOGIC_VECTOR(14 DOWNTO 0) :=(others => '0');
variable DATA_1_n : STD_LOGIC_VECTOR(14 DOWNTO 0) :="101000101000000";

begin
      if (clk'event and clk = '1') then


			DATA_0 <= DATA_0_i;					
			DATA_1 <= DATA_1_i + DATA_0_i;	


			--normalize Data_1 and save amount of shift steps necesarry

			if DATA_0  = "000000000000000" then
				n1_sh <= 0;
				DATA_1_n := "000000000000000";
			elsif (DATA_1(14) = '1') then
				n1_sh <= 0;
				DATA_1_n := DATA_1;
			elsif (DATA_1(13) = '1') then
				n1_sh <= 1;
				DATA_1_n := DATA_1(13 downto 0) & "0";
			elsif (DATA_1(12) = '1') then
				n1_sh <= 2;
				DATA_1_n := DATA_1(12 downto 0) & "00";
			elsif (DATA_1(11) = '1') then
				n1_sh <= 3;
				DATA_1_n := DATA_1(11 downto 0) & "000";
			elsif (DATA_1(10) = '1') then
				n1_sh <= 4;
				DATA_1_n := DATA_1(10 downto 0) & "0000";
			elsif (DATA_1(9) = '1') then
				n1_sh <= 5;
				DATA_1_n := DATA_1(9 downto 0) & "00000";
			elsif(DATA_1(8) = '1') then
				n1_sh <= 6;
				DATA_1_n := DATA_1(8 downto 0) & "000000";
			elsif (DATA_1(7) = '1') then
				n1_sh <= 7;
				DATA_1_n := DATA_1(7 downto 0) & "0000000";
			elsif(DATA_1(6) = '1') then
				n1_sh <= 8;
				DATA_1_n := DATA_1(6 downto 0) & "00000000";
			elsif(DATA_1(5) = '1') then
				n1_sh <= 9;
				DATA_1_n := DATA_1(5 downto 0) & "000000000";
			elsif(DATA_1(4) = '1') then
				n1_sh <= 10;
				DATA_1_n := DATA_1(4 downto 0) & "0000000000";
			elsif(DATA_1(3) = '1') then
				n1_sh <= 11;
				DATA_1_n := DATA_1(3 downto 0) & "00000000000";
			elsif(DATA_1(2) = '1') then
				n1_sh <= 12;
				DATA_1_n := DATA_1(2 downto 0) & "000000000000";
			elsif(DATA_1(1) = '1') then
				n1_sh <= 13;
				DATA_1_n := DATA_1(1 downto 0) & "0000000000000";
			elsif(DATA_1(0) = '1') then
				n1_sh <= 14;
				DATA_1_n := DATA_1(0) & "00000000000000";
			end if;

			--normalize Data_0 and save amount of shift steps necesarry

			if DATA_0  = "000000000000000" then
				n0_sh <= 0;
				DATA_0_n <= "0" & DATA_0;
			elsif (DATA_0(14) = '1') then
				n0_sh <= 0;
				DATA_0_n <= "0" & DATA_0;
			elsif (DATA_0(13) = '1') then
				n0_sh <= 1;
				DATA_0_n <= "0" & DATA_0(13 downto 0) & "0";
			elsif (DATA_0(12) = '1') then
				n0_sh <= 2;
				DATA_0_n <= "0" & DATA_0(12 downto 0) & "00";
			elsif (DATA_0(11) = '1') then
				n0_sh <= 3;
				DATA_0_n <= "0" & DATA_0(11 downto 0) & "000";
			elsif (DATA_0(10) = '1') then
				n0_sh <= 4;
				DATA_0_n <= "0" & DATA_0(10 downto 0) & "0000";
			elsif (DATA_0(9) = '1') then
				n0_sh <= 5;
				DATA_0_n <= "0" & DATA_0(9 downto 0) & "00000";
			elsif(DATA_0(8) = '1') then
				n0_sh <= 6;
				DATA_0_n <= "0" & DATA_0(8 downto 0) & "000000";
			elsif (DATA_0(7) = '1') then
				n0_sh <= 7;
				DATA_0_n <= "0" & DATA_0(7 downto 0) & "0000000";
			elsif(DATA_0(6) = '1') then
				n0_sh <= 8;
				DATA_0_n <= "0" & DATA_0(6 downto 0) & "00000000";
			elsif(DATA_0(5) = '1') then
				n0_sh <= 9;
				DATA_0_n <= "0" & DATA_0(5 downto 0) & "000000000";
			elsif(DATA_0(4) = '1') then
				n0_sh <= 10;
				DATA_0_n <= "0" & DATA_0(4 downto 0) & "0000000000";
			elsif(DATA_0(3) = '1') then
				n0_sh <= 11;
				DATA_0_n <= "0" & DATA_0(3 downto 0) & "00000000000";
			elsif(DATA_0(2) = '1') then
				n0_sh <= 12;
				DATA_0_n <= "0" & DATA_0(2 downto 0) & "000000000000";
			elsif(DATA_0(1) = '1') then
				n0_sh <= 13;
				DATA_0_n <= "0" & DATA_0(1 downto 0) & "0000000000000";
			elsif(DATA_0(0) = '1') then
				n0_sh <= 14;
				DATA_0_n <= "0" & DATA_0(0) & "00000000000000";
			end if;


			DATA_1_h := "0" & DATA_1_n(14 downto 7) & "0000000"; --save upper 8 bits +sign bit in 15 bit vector
			DATA_1_l := "00000000" & DATA_1_n(6 downto 0);		 --save lower 7 bit  +sign bit in 15 bit vector
			adr <="00" & DATA_1_n(14 downto 7);					 --set adresse for the lookup table
			DATA_1_hml <= DATA_1_h - DATA_1_l;						 --get difference of upper and lower bits, DATA_1_hml gets multiplied by DATA_0_n 


			n01_sh <= n0_sh-n1_sh;										 --get difference of shift steps necesarry to normalize denominator and divisor, n0 and n1 max shoulde be 11 => max=11, min=-11
			-- memDO <= BRAM(adr)
			-- multi1 <= DSP(DATA_1_hml * DATA_0_n)


			n01_sh_del <= n01_sh;										 --delay difference of shifts
			mult1_sh <= mult1(31 downto 15); 						 --save 14 bit result of DATA_1_hml * DATA_0_n (not 12 + 1SignBit because of possible error correction), gets multiplied by DATA_1_h_rs 
			DATA_1_h_rs<= "01" & memDO(15 downto 0);            --receive normalized reciproc square of DATA_1 from lookup, 0 is sign, 1 is not saved - normalization
			n_sh <= conv_integer(memDO(21 downto 16));          --receive shift steps of normalized reciproc square from lookup, max should be 24, min = 12


			shift_end <=n01_sh_del+ n_sh+1;                     --add all shift steps, max shoulde be 36 min=1
			-- solution_us <= DSP(mult1_sh * DATA_1_h_rs)

			
			solution_us_del <=solution_us;                      --delay, due to timing constraints in full design
			shift_end_del <= shift_end;								 --delay, due to timing constraints in full design


			test:="000000000" & solution_us_del;					 --9 zeros +1 sign zero, precision 10 bit
			if shift_end_del/=1 then
				adrB <= test(shift_end_del-3 downto shift_end_del-12);--use shifts to get result
			else
				adrB <="0000000000";
			end if;

			result<=memDO_B(31 downto 22);
		
		end if;

end process;

   MULT_MACRO_inst : MULT_MACRO
   generic map (
      DEVICE => "VIRTEX5",    -- Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6" 
      LATENCY => 1,           -- Desired clock cycle latency, 0-4
		WIDTH_A => 16,          -- Multiplier A-input bus width, 1-25 
      WIDTH_B => 16)          -- Multiplier B-input bus width, 1-18
   port map (
      P => mult1,     -- Multiplier ouput bus, width determined by WIDTH_P generic 
      A => DATA_1_hml,     -- Multiplier input A bus, width determined by WIDTH_A generic 
      B => Data_0_n,     -- Multiplier input B bus, width determined by WIDTH_B generic 
      CE => '1',   -- 1-bit active high input clock enable
      CLK => clk, -- 1-bit positive edge clock input
      RST => '0'  -- 1-bit input active high reset
   );

   MULT_MACRO_inst_1 : MULT_MACRO
   generic map (
      DEVICE => "VIRTEX5",    -- Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6" 
      LATENCY => 1,           -- Desired clock cycle latency, 0-4
		WIDTH_A =>17,          -- Multiplier A-input bus width, 1-25 
      WIDTH_B => 18)          -- Multiplier B-input bus width, 1-18
   port map (
      P => solution_us,     -- Multiplier ouput bus, width determined by WIDTH_P generic 
      A => mult1_sh,     -- Multiplier input A bus, width determined by WIDTH_A generic 
      B => DATA_1_h_rs,     -- Multiplier input B bus, width determined by WIDTH_B generic 
      CE => '1',   -- 1-bit active high input clock enable
      CLK => clk, -- 1-bit positive edge clock input
      RST => '0'  -- 1-bit input active high reset
   );


   BRAM_TDP_MACRO_inst : BRAM_TDP_MACRO
   generic map (
      BRAM_SIZE => "36Kb", -- Target BRAM, "18Kb" or "36Kb" 
      DEVICE => "VIRTEX5", -- Target Device: "VIRTEX5", "VIRTEX6", "SPARTAN6" 
      DOA_REG => 0, -- Optional port A output register (0 or 1)
      DOB_REG => 0, -- Optional port B output register (0 or 1)
      INIT_A => X"ABCDEFF12", -- Initial values on A output port
      INIT_B => X"ABCDEFF12", -- Initial values on B output port
      INIT_FILE => "NONE",
      READ_WIDTH_A => 36,   -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
      READ_WIDTH_B => 36,   -- Valid values are 1-36 (19-36 only valid when BRAM_SIZE="36Kb")
      SIM_COLLISION_CHECK => "ALL", -- Collision check enable "ALL", "WARNING_ONLY", 
                                    -- "GENERATE_X_ONLY" or "NONE" 
      SIM_MODE => "FAST", -- Simulation: "SAFE" vs "FAST",                                  -- era SAFE
                          -- see "Synthesis and Simulation Design Guide" for details
      SRVAL_A => X"000000000",   -- Set/Reset value for A port output
      SRVAL_B => X"000000000",   -- Set/Reset value for B port output
      WRITE_MODE_A => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE" 
      WRITE_MODE_B => "WRITE_FIRST", -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE" 
      WRITE_WIDTH_A => 36, -- Valid values are 1, 2, 4, 9, 18 or 36 (36 only valid when BRAM_SIZE="36Kb")
      WRITE_WIDTH_B => 36, -- Valid values are 1, 2, 4, 9, 18 or 36 (36 only valid when BRAM_SIZE="36Kb")
      -- The following INIT_xx declarations specify the initial contents of the RAM

		INIT_00 => b"0000000111010110010011100101111000000001100101101100011100011100000000010101010101000111101011100000000100010100000000000000000000000000110101001100011100011100000000001001001000000000000000000000000001010000000000000000000000000000000000000000000000000000",
		INIT_01 => b"0000001111011000001000110100010100000011100110000100111001011110000000110101100010000011110010010000001100011000110001110001110000000010110101110000111011001111000000101001011101000111101011100000001001010111100101001000101100000010000101100000000000000000",
		INIT_02 => b"0000010111011010111011111000101100000101100110010000111011001111000001010101100100101001001101110000010100011001010001111010111000000100110110010110101100010100000001001001100110010100100010110000010001011001110001011000100100000100000110000000000000000000",
		INIT_03 => b"0000011111011010000100001100100000000111100110100010001101000101000001110101101000110111101101000000011100011010010011100101111000000110110110100110011110011000000001101001101010000011110010010000011001011010101000110110111000000110000110101100011100011100",
		INIT_04 => b"0000100111011011010110001011001100001001100110110110101100010100000010010101101101111110111110000000100100011011100101001000101100001000110110111010101111111101000010001001101111000101100010010000100001011011111000010111000000001000000110100000000000000000",
		INIT_05 => b"0000101111011100110110101010111000001011100111001110111110001011000010110101101100000010111010000000101100011011000011101100111100001010110110110001101110001101000010101001101100101001001101110000101001011011001101111110001100001010000110110100011110101110",
		INIT_06 => b"0000110111011100010110101010001000001101100111000110011110011000000011010101110001110101010010100000110100011100100000111100100100001100110111001001001100100100000011001001110010100011011011100000110001011100101101001011100100001100000111001100011100011100",
		INIT_07 => b"0000111111011100000010000011000100001111100111000001000011001000000011110101110000011001110011000000111100011100001000110100010100001110110111000010110100111010000011101001110000110111101101000000111001011100010000101011110000001110000111000100111001011110",
		INIT_08 => b"0001000111011101101000000000010000010001100111011010101111111101000100010101110110111000011111000001000100011101110001011000100100010000110111011101001100101100000100001001110111100001011100000001000001011101111100000101111000010000000111000000000000000000",
		INIT_09 => b"0001001111011101010100000000011100010011100111010101100010110011000100110101110101100001101101010001001100011101011010110001010000010010110111010111010011010011000100101001110101111110111110000001001001011101100010011000100100010010000111011001010010001011",
		INIT_0a => b"0001010111011101000101010001001000010101100111010001101110001101000101010101110100100010010000110001010100011101001010010011011100010100110111010011000001101011000101001001110100110111111000110001010001011101001111111010001100010100000111010100011110101110",
		INIT_0b => b"0001011111011110110100001011111000010111100111101101101010101110000101110101111011100100111100100001011100011110111011111000101100010110110111101111101001111111000101101001110100000010111010000001011001011101000010001100001000010110000111010000111011001111",
		INIT_0c => b"0001100111011110100010110101101000011001100111101001001100100100000110010101111010011011001010100001100100011110101000110110111000011000110111101010101111110010000110001001111010110100101110010001100001011110101111011100011000011000000111101100011100011100",
		INIT_0d => b"0001101111011110010101000110101100011011100111100101101010100010000110110101111001100001000001100001101100011110011001111001100000011010110111100110111001011000000110101001111001110101010010100001101001011110011111000110111100011010000111101000001111001001",
		INIT_0e => b"0001110111011110001010000010111100011101100111100010110100111010000111010101111000110010011001100001110100011110001101111011010000011100110111100011110100100110000111001001111001000010101111000001110001011110010010000111100100011100000111100100111001011110",
		INIT_0f => b"0001111111011110000001000000110000011111100111100000100000110001000111110101111000001100011011110001111100011110000100001100100000011110110111100001010100111100000111101001111000011001110011000001111001011110000111100111101000011110000111100010001101000101",
		INIT_10 => b"0010000111011111110011000100011100100001100111111101001100101100001000010101111111011010001110100010000100011111111000010111000000100000110111111110100011010001001000001001111111110000010111100010000001011111111110000001011100100000000111100000000000000000",
		INIT_11 => b"0010001111011111100110100011100000100011100111111010000000000100001000110101111110100101111100000010001100011111101010111111110100100010110111111011001000101011001000101001111110111000011111000010001001011111101111101111000000100010000111111100010110001001",
		INIT_12 => b"0010010111011111011011111110011100100101100111110111010011010011001001010101111101111001110110010010010100011111011111101111100000100100110111111000010000110011001001001001111110001001100010010010010001011111100011101111101100100100000111111001010010001011",
		INIT_13 => b"0010011111011111010010111101000000100111100111110101000000000111001001110101111101010100010100100010011100011111010110001011001100100110110111110101110100101001001001101001111101100001101101010010011001011111011001100101100100100110000111110110101100010100",
		INIT_14 => b"0010100111011111001011001100100100101001100111110011000001101011001010010101111100110100000111110010100100011111001101111110001100101000110111110011101110111010001010001001111100111111101000110010100001011111010000111001111100101000000111110100011110101110",
		INIT_15 => b"0010101111011111000100011110100100101011100111110001010100010010001010110101111100011000010010000010101100011111000110111000110100101010110111110001111011100000001010101001111100100010010000110010101001011111001001011011010100101010000111110010100100110111",
		INIT_16 => b"0010110111100000111101001111101000101101101000001111101001111111001011010101111100000000000011100010110100011111000000101110100000101100110111110000010111001110001011001001111100001000110000100010110001011111000010111100001000101100000111110000111011001111",
		INIT_17 => b"0010111111100000110010111110001100101111101000001101000010111110001011110110000011010101101011000010111100100000110110101010111000101110111000001101111111000110001011101010000011100100111100100010111001100000111010100011010000101110001000001110111110001011",
		INIT_18 => b"0011000111100000101001111010100000110001101000001010101111110010001100010110000010110000010011010011000100100000101101001011100100110000111000001011100100110111001100001010000010111101110001100011000001100000110000100110100000110000001000001100011100011100",
		INIT_19 => b"0011001111100000100001111000101000110011101000001000101101011010001100110110000010001111001110000011001100100000100100110010010000110010111000001001011100100000001100101010000010011011001010100011001001100000100111110100010000110010001000001010001101101110",
		INIT_1a => b"0011010111100000011010101111001000110101101000000110111001011000001101010110000001110001110010110011010100100000011101010100101000110100111000000111100011010110001101001010000001111100011011110011010001100000100000000001010100110100001000001000001111001001",
		INIT_1b => b"0011011111100000010100010101111100110111101000000101010001101011001101110110000001010111100000010011011100100000010110101010001000110110111000000101110111001111001101101010000001100001000001100011011001100000011001000100100100110110001000000110011110011000",
		INIT_1c => b"0011100111100000001110100110100000111001101000000011110100100110001110010110000000111111111011000011100100100000010000101011110000111000111000000100010110010110001110001010000001001000011110010011100001100000010010110110011000111000001000000100111001011110",
		INIT_1d => b"0011101111100000001001011011011000111011101000000010100000101111001110110110000000101010101100010011101100100000001011010011101000111010111000000010111111001100001110101010000000110010011001100011101001100000001101010000100100111010001000000011011110110100",
		INIT_1e => b"0011110111100000000100101111111000111101101000000001010100111100001111010110000000010111100000000011110100100000000110011100110000111100111000000001110000011111001111001010000000011110011110100011110001100000001000001101101100111100001000000010001101000101",
		INIT_1f => b"0011111111100000000000100000001100111111101000000000010000001100001111110110000000000110000110110011111100100000000010000011000100111110111000000000101001001101001111101010000000001100011011110011111001100000000011101001100000111110001000000001000011001000",
		INIT_20 => b"0100000111100001111001010001101101000001101000011110100011010001010000010110000111101100100100100100000100100001111100000101111001000000111000011111010000110101010000001010000111111000000101110100000001100001111111000000010101000000001000000000000000000000",
		INIT_21 => b"0100001111100001110010001110001101000011101000011100110001000111010000110110000111001111101101010100001100100001110100110010110001000010111000011101011010101110010000101010000111011010001110100100001001100001110111011101000001000010001000011110000101110000",
		INIT_22 => b"0100010111100001101011110001000001000101101000011011001000101011010001010110000110110101010011110100010100100001101110000111110001000100111000011011101110110001010001001010000110111110111100000100010001100001110000100011100001000100001000011100010110001001",
		INIT_23 => b"0100011111100001100101110101111001000111101000011001101000111000010001110110000110011101000110100100011100100001101000000000010001000110111000011010001011110110010001101010000110100101111100000100011001100001101010001111001101000110001000011010101111111101",
		INIT_24 => b"0100100111100001100000011001001001001001101000011000010000110011010010010110000110000110110110100100100100100001100010011000100101001000111000011000110000111110010010001010000110001110111110110100100001100001100100011011111101001000001000011001010010001011",
		INIT_25 => b"0100101111100001011011010111101101001011101000010110111111100111010010110110000101110010010110100100101100100001011101001101001101001010111000010111011101010011010010101010000101111001110110010100101001100001011111000110010101001010001000010111111011111000",
		INIT_26 => b"0100110111100001010110101110101101001101101000010101110100101001010011010110000101011111011011000100110100100001011000011011010101001100111000010110010000000100010011001010000101100110010110010100110001100001011010001011010001001100001000010110101100010100",
		INIT_27 => b"0100111111100001010010011011110001001111101000010100101111010000010011110110000101001101111010010100111100100001010100000000011101001110111000010101001000101010010011101010000101010100010100100100111001100001010101101000000001001110001000010101100010110011",
		INIT_28 => b"0101000111100001001110011100110101010001101000010011101110111010010100010110000100111101101011000101000100100001001111111010001101010000111000010100000110011111010100001010000101000011100111110101000001100001010001011010010001010000001000010100011110101110",
		INIT_29 => b"0101001111100001001010101111111001010011101000010010110011001001010100110110000100101110100110000101001100100001001100000110101101010010111000010011001001000011010100101010000100110100000111110101001001100001001101011111111101010010001000010011011111100011",
		INIT_2a => b"0101010111100001000111010011010101010101101000010001111011100000010101010110000100100000100100000101010100100001001000100100001101010100111000010010001111111010010101001010000100100101101101010101010001100001001001110111010001010100001000010010100100110111",
		INIT_2b => b"0101011111100001000100000101101001010111101000010001000111101001010101110110000100010011011111000101011100100001000101010001001001010110111000010001011010101011010101101010000100011000010010000101011001100001000110011110100101010110001000010001101110001101",
		INIT_2c => b"0101100111100001000001000101101001011001101000010000010111001110010110010110000100000111010001100101100100100001000010001100001001011000111000010000101001000000010110001010000100001011110000100101100001100001000011010100011101011000001000010000111011001111",
		INIT_2d => b"0101101111100010111100100100000001011011101000101111010011111010010110110110001011110111101110010101101100100010111110100111111101011010111000101111110101001010010110101010000100000000000011100101101001100001000000010111100101011010001000010000001011101000",
		INIT_2e => b"0101110111100010110111010011011101011101101000101101111111000110010111010110001011100010010110010101110100100010111001001111001001011100111000101110011110010000010111001010001011101010001101000101110001100010111011001101110101011100001000101110111110001011",
		INIT_2f => b"0101111111100010110010010111110101011111101000101100101111100011010111110110001011001110010011100101111100100010110100001011111001011110111000101101001100110010010111101010001011010101101011000101111001100010110110000010101101011110001000101101101010101110",
		INIT_30 => b"0110000111100010101101101111011001100001101000101011100100110111011000010110001010111011011111000110000100100010101111011100011001100000111000101100000000010101011000001010001011000010011010000110000001100010110001001011111101100000001000101100011100011100",
		INIT_31 => b"0110001111100010101001011000100101100011101000101010011110101000011000110110001010101001110010110110001100100010101010111111001001100010111000101010111000011101011000101010001010110000010011010110001001100010101100101000000101100010001000101011010010111001",
		INIT_32 => b"0110010111100010100101010010000001100101101000101001011100100000011001010110001010011001001000110110010100100010100110110010101001100100111000101001110100110101011001001010001010011111010001000110010001100010101000010101011101100100001000101010001101101110",
		INIT_33 => b"0110011111100010100001011010100001100111101000101000011110001010011001110110001010001001011100000110011100100010100010110101101001100110111000101000110101000111011001101010001010001111001110000110011001100010100100010010110001100110001000101001001100100100",
		INIT_34 => b"0110100111100010011101110000111101101001101000100111100011010110011010010110001001111010101000010110100100100010011111000110111101101000111000100111111001000000011010001010001010000000000101010110100001100010100000011110110101101000001000101000001111001001",
		INIT_35 => b"0110101111100010011010010100001101101011101000100110101011110010011010110110001001101100101001000110101100100010011011100101100001101010111000100111000000010000011010101010001001110001110010110110101001100010011100111000100101101010001000100111010101001010",
		INIT_36 => b"0110110111100010010111000011011101101101101000100101110111001111011011010110001001011111011010010110110100100010011000010000011001101100111000100110001010100110011011001010001001100100010010010110110001100010011001011110111101101100001000100110011110011000",
		INIT_37 => b"0110111111100010010011111101110101101111101000100101000101011111011011110110001001010010111001000110111100100010010101000110101101101110111000100101010111110101011011101010001001010111100000010110111001100010010110010001000101101110001000100101101010100010",
		INIT_38 => b"0111000111100010010001000010100001110001101000100100010110010110011100010110001001000111000001100111000100100010010010000111100101110000111000100100100111101111011100001010001001001011011001100111000001100010010011001110000101110000001000100100111001011110",
		INIT_39 => b"0111001111100010001110010000110101110011101000100011101001101000011100110110001000111011110001100111001100100010001111010010011001110010111000100011111010001000011100101010001000111111111011000111001001100010010000010101001101110010001000100100001010111100",
		INIT_3a => b"0111010111100010001011101000001001110101101000100010111111001100011101010110001000110001000110000111010100100010001100100110011001110100111000100011001110110110011101001010001000110101000010010111010001100010001101100101110101110100001000100011011110110100",
		INIT_3b => b"0111011111100010001001000111110101110111101000100010010110110110011101110110001000100110111100100111011100100010001010000010111101110110111000100010100101101111011101101010001000101010101100010111011001100010001010111111010001110110001000100010110100111010",
		INIT_3c => b"0111100111100010000110101111010101111001101000100001110000011111011110010110001000011101010010110111100100100010000111100111101001111000111000100001111110101010011110001010001000100000110110110111100001100010001000100000111101111000001000100010001101000101",
		INIT_3d => b"0111101111100010000100011110001001111011101000100001001011111110011110110110001000010100000111000111101100100010000101010011110001111010111000100001011001011101011110101010001000010111100000000111101001100010000110001010010101111010001000100001100111001100",
		INIT_3e => b"0111110111100010000010010011111001111101101000100000101001001101011111010110001000001011010111010111110100100010000011000110111101111100111000100000110110000011011111001010001000001110100110000111110001100010000011111010111101111100001000100001000011001000",
		INIT_3f => b"0111111111100010000000010000000001111111101000100000001000000011011111110110001000000011000001100111111100100010000001000000110001111110111000100000010100010010011111101010001000000110000110110111111001100010000001110010010101111110001000100000100000110001",
		INIT_40 => b"1000000111100011111100100100100010000001101000111111010000110101100000010110001111110110001001011000000100100011111110000001011110000000111000111111101000001101100000001010001111111100000001011000000001100011111111100000000110000000001000100000000000000000",
		INIT_41 => b"1000001111100011111000110100010010000011101000111110010100011011100000110110001111100110111101011000001100100011111010001101000110000010111000111110101010110000100000101010001111101100100100101000001001100011111011100111011010000010001000111111000001011110",
		INIT_42 => b"1000010111100011110101001110110010000101101000111101011010101110100001010110001111011000011100111000010100100011110110100011101010000100111000111101110000000011100001001010001111011101110100001000010001100011110111111001111110000100001000111110000101110000",
		INIT_43 => b"1000011111100011110001110011010110000111101000111100100011100011100001110110001111001010100101001000011100100011110011000100011110000110111000111100110111111101100001101010001111001111101101011000011001100011110100010110111110000110001000111101001100101100",
		INIT_44 => b"1000100111100011101110100001010110001001101000111011101110110001100010010110001110111101010100001000100100100011101111101111000010001000111000111100000010010011100010001010001111000010001110001000100001100011110000111101111110001000001000111100010110001001",
		INIT_45 => b"1000101111100011101011011000010110001011101000111010111100010000100010110110001110110000100111001000101100100011101100100010101110001010111000111011001110111100100010101010001110110101010011111000101001100011101101101110010010001010001000111011100001111100",
		INIT_46 => b"1000110111100011101000010111110010001101101000111010001011110110100011010110001110100100011100101000110100100011101001011111000010001100111000111010011101110000100011001010001110101000111100111000110001100011101010100111011110001100001000111010101111111101",
		INIT_47 => b"1000111111100011100101011111001110001111101000111001011101011110100011110110001110011000110010101000111100100011100110100011100010001110111000111001101110101000100011101010001110011101000110101000111001100011100111101000111010001110001000111010000000000100",
		INIT_48 => b"1001000111100011100010101110001110010001101000111000110000111110100100010110001110001101100111001001000100100011100011101111101110010000111000111001000001011100100100001010001110010001101111111001000001100011100100110010010010010000001000111001010010001011",
		INIT_49 => b"1001001111100011100000000100010010010011101000111000000110010010100100110110001110000010111000011001001100100011100001000011001110010010111000111000010110000110100100101010001110000110110110101001001001100011100010000011000110010010001000111000100110001001",
		INIT_4a => b"1001010111100011011101100001001010010101101000110111011101010011100101010110001101111000100101011001010100100011011110011101100110010100111000110111101100011110100101001010001101111100011001011001010001100011011111011010111010010100001000110111111011111000",
		INIT_4b => b"1001011111100011011011000100011110010111101000110110110101111011100101110110001101101110101100001001011100100011011011111110011110010110111000110111000100100000100101101010001101110010010110101001011001100011011100111001011010010110001000110111010011010011",
		INIT_4c => b"1001100111100011011000101101110010011001101000110110010000000100100110010110001101100101001011101001100100100011011001100101100110011000111000110110011110000110100110001010001101101000101101001001100001100011011010011110001110011000001000110110101100010100",
		INIT_4d => b"1001101111100011010110011100111010011011101000110101101011101011100110110110001101011100000010011001101100100011010111010010100110011010111000110101111001001010100110101010001101011111011011001001101001100011011000001001000010011010001000110110000110110101",
		INIT_4e => b"1001110111100011010100010001100010011101101000110101001000101010100111010110001101010011001111011001110100100011010101000101001010011100111000110101010101101000100111001010001101010110100000001001110001100011010101111001100010011100001000110101100010110011",
		INIT_4f => b"1001111111100011010010001011010010011111101000110100100110111100100111110110001101001010110001101001111100100011010010111101000010011110111000110100110011011100100111101010001101001101111010011001111001100011010011101111011110011110001000110101000000000111",
		INIT_50 => b"1010000111100011010000001010000010100001101000110100000110011111101000010110001101000010100111101010000100100011010000111001111110100000111000110100010010100001101000001010001101000101101001001010000001100011010001101010100010100000001000110100011110101110",
		INIT_51 => b"1010001111100011001110001101011110100011101000110011100111001101101000110110001100111010110000111010001100100011001110111011101010100010111000110011110010110011101000101010001100111101101011001010001001100011001111101010011110100010001000110011111110100011",
		INIT_52 => b"1010010111100011001100010101011010100101101000110011001001000011101001010110001100110011001100001010010100100011001101000001111110100100111000110011010100001110101001001010001100110101111111111010010001100011001101101111000110100100001000110011011111100011",
		INIT_53 => b"1010011111100011001010100001101010100111101000110010101011111110101001110110001100101011111000111010011100100011001011001100100110100110111000110010110110110000101001101010001100101110100110001010011001100011001011111000000110100110001000110011000001101011",
		INIT_54 => b"1010100111100011001000110001111010101001101000110010001111111010101010010110001100100100110101111010100100100011001001011011010110101000111000110010011010010100101010001010001100100111011101001010100001100011001010000101010110101000001000110010100100110111",
		INIT_55 => b"1010101111100011000111000110000010101011101000110001110100110101101010110110001100011110000010101010101100100011000111101110000010101010111000110001111110111000101010101010001100100000100100001010101001100011001000010110100110101010001000110010001001000011",
		INIT_56 => b"1010110111100011000101011101111010101101101000110001011010101011101011010110001100010111011110011010110100100011000110000100100010101100111000110001100100011000101011001010001100011001111010011010110001100011000110101011101010101100001000110001101110001101",
		INIT_57 => b"1010111111100011000011111001010010101111101000110001000001011010101011110110001100010001001000011010111100100011000100011110100110101110111000110001001010110010101011101010001100010011011111001010111001100011000101000100011010101110001000110001010100010010",
		INIT_58 => b"1011000111100011000010011000000010110001101000110000101001000000101100010110001100001011000000001011000100100011000010111100001010110000111000110000110010000100101100001010001100001101010001111011000001100011000011100000101010110000001000110000111011001111",
		INIT_59 => b"1011001111100011000000111010000010110011101000110000010001011010101100110110001100000101000101001011001100100011000001011100111010110010111000110000011010001010101100101010001100000111010001101011001001100011000010000000010010110010001000110000100011000010",
		INIT_5a => b"1011010111100100111110111110010010110101101001001111110101001010101101010110010011111110101100101011010100100011000000000000111010110100111000110000000011000011101101001010001100000001011110011011010001100011000000100011000010110100001000110000001011101000",
		INIT_5b => b"1011011111100100111100001110010110110111101001001111001001000000101101110110010011110011100111001011011100100100111101001111101010110110111001001111011001011001101101101010010011110111101110011011011001100100111110010001101110110110001001001111101001111111",
		INIT_5c => b"1011100111100100111001100100000010111001101001001110011110010000101110010110010011101000111000011011100100100100111010100011010010111000111001001110101110000111101110001010010011101100110111011011100001100100111011100011001110111000001001001110111110001011",
		INIT_5d => b"1011101111100100110110111111001010111011101001001101110100110111101110110110010011011110011111101011101100100100110111111100011010111010111001001110000100001111101110101010010011100010010110011011101001100100111000111010010110111010001001001110010011110010",
		INIT_5e => b"1011110111100100110100011111011110111101101001001101001100110010101111010110010011010100011011111011110100100100110101011010110010111100111001001101011011101011101111001010010011011000001010111011110001100100110110010110110010111100001001001101101010101110",
		INIT_5f => b"1011111111100100110010000100110010111111101001001100100101111101101111110110010011001010101100001011111100100100110010111110001110111110111001001100110100011000101111101010010011001110010011101011111001100100110011111000010110111110001001001101000010111110",
		INIT_60 => b"1100000111100100101111101110110111000001101001001100000000010101110000010110010011000001001111101100000100100100110000100110100011000000111001001100001110010011110000001010010011000100101111111100000001100100110001011110110111000000001001001100011100011100",
		INIT_61 => b"1100001111100100101101011101011111000011101001001011011011110110110000110110010010111000000101101100001100100100101110010011011111000010111001001011101001011001110000101010010010111011011111001100001001100100101111001010000111000010001001001011110111000110",
		INIT_62 => b"1100010111100100101011010000011111000101101001001010111000011101110001010110010010101111001101011100010100100100101100000100110111000100111001001011000101100110110001001010010010110010100000011100010001100100101100111001110011000100001001001011010010111001",
		INIT_63 => b"1100011111100100101001000111101111000111101001001010010110001001110001110110010010100110100110001100011100100100101001111010100011000110111001001010100010111001110001101010010010101001110010111100011001100100101010101101111011000110001001001010101111110010",
		INIT_64 => b"1100100111100100100111000010111111001001101001001001110100110101110010010110010010011110001111001100100100100100100111110100010011001000111001001010000001001101110010001010010010100001010101111100100001100100101000100110001011001000001001001010001101101110",
		INIT_65 => b"1100101111100100100101000010001011001011101001001001010100100000110010110110010010010110000111111100101100100100100101110010000011001010111001001001100000100001110010101010010010011001001000111100101001100100100110100010011011001010001001001001101100101010",
		INIT_66 => b"1100110111100100100011000101000011001101101001001000110101000111110011010110010010001110001111111100110100100100100011110011100011001100111001001001000000110010110011001010010010010001001011001100110001100100100100100010100011001100001001001001001100100100",
		INIT_67 => b"1100111111100100100001001011100011001111101001001000010110101000110011110110010010000110100110011100111100100100100001111000101011001110111001001000100001111101110011101010010010001001011100001100111001100100100010100110010111001110001001001000101101011010",
		INIT_68 => b"1101000111100100011111010101011111010001101001000111111001000000110100010110010001111111001010101101000100100100100000000001010111010000111001001000000100000001110100001010010010000001111011011101000001100100100000101101101111010000001001001000001111001001",
		INIT_69 => b"1101001111100100011101100010110011010011101001000111011100001111110100110110010001110111111100101101001100100100011110001101011011010010111001000111100110111011110100101010010001111010101000011101001001100100011110111000100011010010001001000111110001101111",
		INIT_6a => b"1101010111100100011011110011010011010101101001000111000000010000110101010110010001110000111011011101010100100100011100011100101111010100111001000111001010101010110101001010010001110011100010011101010001100100011101000110100111010100001001000111010101001010",
		INIT_6b => b"1101011111100100011010000110110111010111101001000110100101000011110101110110010001101010000110101101011100100100011010101111001011010110111001000110101111001010110101101010010001101100101001001101011001100100011011010111111011010110001001000110111001011000",
		INIT_6c => b"1101100111100100011000011101011011011001101001000110001010100110110110010110010001100011011101111101100100100100011001000100100111011000111001000110010100011100110110001010010001100101111011111101100001100100011001101100001111011000001001000110011110011000",
		INIT_6d => b"1101101111100100010110110110110111011011101001000101110000110111110110110110010001011101000000111101101100100100010111011100111111011010111001000101111010011100110110101010010001011111011010011101101001100100011000000011011111011010001001000110000100000110",
		INIT_6e => b"1101110111100100010101010010111111011101101001000101010111110101110111010110010001010110101110111101110100100100010101111000000111011100111001000101100001001001110111001010010001011001000100011101110001100100010110011101100111011100001001000101101010100010",
		INIT_6f => b"1101111111100100010011110001110111011111101001000100111111011101110111110110010001010000100111101101111100100100010100010101111111011110111001000101001000100001110111101010010001010010111001001101111001100100010100111010011111011110001001000101010001101011",
		INIT_70 => b"1110000111100100010010010011010011100001101001000100100111101111111000010110010001001010101010101110000100100100010010110110011011100000111001000100110000100011111000001010010001001100111000011110000001100100010011011001111111100000001001000100111001011110",
		INIT_71 => b"1110001111100100010000110111001011100011101001000100010000101000111000110110010001000100110111111110001100100100010001011001011011100010111001000100011001001110111000101010010001000111000001101110001001100100010001111100000011100010001001000100100001111001",
		INIT_72 => b"1110010111100100001111011101011111100101101001000011111010001000111001010110010000111111001110101110010100100100001111111110110011100100111001000100000010100000111001001010010001000001010100111110010001100100010000100000100011100100001001000100001010111100",
		INIT_73 => b"1110011111100100001110000110000011100111101001000011100100001101111001110110010000111001101110101110011100100100001110100110100011100110111001000011101100010111111001101010010000111011110001101110011001100100001111000111011011100110001001000011110100100110",
		INIT_74 => b"1110100111100100001100110000111011101001101001000011001110110110111010010110010000110100010111111110100100100100001101010000100111101000111001000011010110110011111010001010010000110110010111011110100001100100001101110000100011101000001001000011011110110100",
		INIT_75 => b"1110101111100100001011011101111011101011101001000010111010000010111010110110010000101111001001101110101100100100001011111100110011101010111001000011000001110001111010101010010000110001000110001110101001100100001100011011111011101010001001000011001001100110",
		INIT_76 => b"1110110111100100001010001100111111101101101001000010100101101111111011010110010000101010000100001110110100100100001010101011000111101100111001000010101101010010111011001010010000101011111101001110110001100100001011001001011111101100001001000010110100111010",
		INIT_77 => b"1110111111100100001000111110000011101111101001000010010001111101111011110110010000100101000110011110111100100100001001011011011011101110111001000010011001010100111011101010010000100110111100101110111001100100001001111001000011101110001001000010100000101111",
		INIT_78 => b"1111000111100100000111110001000111110001101001000001111110101010111100010110010000100000010000101111000100100100001000001101101111110000111001000010000101110101111100001010010000100010000011111111000001100100001000101010101011110000001001000010001101000101",
		INIT_79 => b"1111001111100100000110100110000011110011101001000001101011110101111100110110010000011011100010101111001100100100000111000001111111110010111001000001110010110101111100101010010000011101010010111111001001100100000111011110001011110010001001000001111001111010",
		INIT_7a => b"1111010111100100000101011100110011110101101001000001011001011101111101010110010000010110111011111111010100100100000101111000000011110100111001000001100000010011111101001010010000011000101001011111010001100100000110010011100111110100001001000001100111001100",
		INIT_7b => b"1111011111100100000100010101010111110111101001000001000111100010111101110110010000010010011100001111011100100100000100101111111011110110111001000001001110001101111101101010010000010100000111001111011001100100000101001010110011110110001001000001010100111100",
		INIT_7c => b"1111100111100100000011001111100111111001101001000000110110000011111110010110010000001110000011011111100100100100000011101001100011111000111001000000111100100011111110001010010000001111101011111111100001100100000100000011101111111000001001000001000011001000",
		INIT_7d => b"1111101111100100000010001011011111111011101001000000100100111110111110110110010000001001110001011111101100100100000010100100110111111010111001000000101011010101111110101010010000001011010111011111101001100100000010111110011011111010001001000000110001101111",
		INIT_7e => b"1111110111100100000001001000111111111101101001000000010100010010111111010110010000000101100101111111110100100100000001100001101111111100111001000000011010100000111111001010010000000111001001011111110001100100000001111010101111111100001001000000100000110001",
        INIT_7f => b"1111111111100100000000001000000011111111101001000000000100000000111111110110010000000001100000011111111100100100000000100000001111111110111001000000001010000100111111101010010000000011000001101111111001100100000000111000100111111110001001000000010000001100",

      
      -- The next set of INITP_xx are for the parity bits
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      
      -- The next set of INIT_xx are valid when configured as 36Kb
      INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000")
    port map (
      DOA => memDO,       -- Output port-A data
      DOB => memDO_B,       -- Output port-B data
      ADDRA =>adr,   -- Input port-A address
      ADDRB => adrB,   -- Input port-B address
      CLKA => clk,     -- Input port-A clock
      CLKB => clk,     -- Input port-B clock
      DIA => test2,       -- Input port-A data
      DIB => test2,       -- Input port-B data
      ENA => '1',       -- Input port-A enable
      ENB => '1' ,     -- Input port-B enable
      REGCEA =>'0', -- Input port-A output register enable
      REGCEB => '0',-- Input port-B output register enable
      RSTA =>'0',     -- Input port-A reset
      RSTB =>'0',     -- Input port-B reset
      WEA => test3,       -- Input port-A write enable
      WEB => test3        -- Input port-B write enable
   );


--  port map (
--    DO => memDO,      -- Output data
--    ADDR => adr,  -- Input address
--    CLK => 	clk,    -- Input clock
--    DI => 	test2,      -- Input data port  
--    EN =>	'1',      -- Input RAM enable
--    REGCE => '0', -- Input output register enable
--    RST => '0',    -- Input reset
--    WE => test3       -- Input write enable
-- );

			
end Behavioral;
