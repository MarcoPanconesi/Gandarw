------------------------------------------------------------------------------
--$Date: 2010/06/25 15:58:07 $
--$Revision: 1.7 $
------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /
-- \   \   \/     Vendor : Xilinx
--  \   \         Version : 2.1
--  /   /         Application : RocketIO GTP Transceiver Wizard
-- /___/   /\     Filename : single_channel_aurora_xc5vsx95t_top.vhd
-- \   \  /  \
--  \___\/\___\
--
--
-- Module SINGLE_CHANNEL_AURORA_XC5VSX95T_TOP
-- Generated by Xilinx RocketIO GTP Transceiver Wizard
-- 
-- 
-- (c) Copyright 2006-2010 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;


--***********************************Entity Declaration************************

entity SINGLE_CHANNEL_AURORA_XC5VSX95T_TOP is
generic
(
    EXAMPLE_CONFIG_INDEPENDENT_LANES        : integer   := 1;
    EXAMPLE_LANE_WITH_START_CHAR            : integer   := 0;
    EXAMPLE_WORDS_IN_BRAM                   : integer   := 512;
    EXAMPLE_SIM_MODE                        : string    := "FAST";
    EXAMPLE_SIM_GTPRESET_SPEEDUP            : integer   := 1;
    EXAMPLE_SIM_PLL_PERDIV2                 : bit_vector:= x"141";
    EXAMPLE_USE_CHIPSCOPE                   : integer   := 1     -- Set to 1 to use Chipscope to drive resets
);
port
(
    TILE0_REFCLK_PAD_N_IN                   : in   std_logic;
    TILE0_REFCLK_PAD_P_IN                   : in   std_logic;
    GTPRESET_IN                             : in   std_logic;
    TILE0_PLLLKDET_OUT                      : out  std_logic;
    TRACK_DATA_OUT                          : out  std_logic;
    RXN_IN                                  : in   std_logic_vector(1 downto 0);
    RXP_IN                                  : in   std_logic_vector(1 downto 0);
    TXN_OUT                                 : out  std_logic_vector(1 downto 0);
    TXP_OUT                                 : out  std_logic_vector(1 downto 0)
    
);

    attribute X_CORE_INFO : string;
    attribute X_CORE_INFO of SINGLE_CHANNEL_AURORA_XC5VSX95T_TOP : entity is "v5_gtpwizard_v2_1, Coregen v12.1";

end SINGLE_CHANNEL_AURORA_XC5VSX95T_TOP;
    
architecture RTL of SINGLE_CHANNEL_AURORA_XC5VSX95T_TOP is

--**************************Component Declarations*****************************


component SINGLE_CHANNEL_AURORA_XC5VSX95T 
generic
(
    -- Simulation attributes
    WRAPPER_SIM_MODE                : string    := "FAST"; -- Set to Fast Functional Simulation Model    
    WRAPPER_SIM_GTPRESET_SPEEDUP    : integer   := 0; -- Set to 1 to speed up sim reset
    WRAPPER_SIM_PLL_PERDIV2         : bit_vector:= x"141" -- Set to the VCO Unit Interval time
);
port
(
    
    --_________________________________________________________________________
    --_________________________________________________________________________
    --TILE0  (Location)

    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    TILE0_RXCHARISCOMMA0_OUT                : out  std_logic_vector(1 downto 0);
    TILE0_RXCHARISCOMMA1_OUT                : out  std_logic_vector(1 downto 0);
    TILE0_RXCHARISK0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXCHARISK1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXDISPERR0_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXDISPERR1_OUT                    : out  std_logic_vector(1 downto 0);
    TILE0_RXNOTINTABLE0_OUT                 : out  std_logic_vector(1 downto 0);
    TILE0_RXNOTINTABLE1_OUT                 : out  std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    TILE0_RXBYTEISALIGNED0_OUT              : out  std_logic;
    TILE0_RXBYTEISALIGNED1_OUT              : out  std_logic;
    TILE0_RXENMCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENMCOMMAALIGN1_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN0_IN               : in   std_logic;
    TILE0_RXENPCOMMAALIGN1_IN               : in   std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    TILE0_RXDATA0_OUT                       : out  std_logic_vector(15 downto 0);
    TILE0_RXDATA1_OUT                       : out  std_logic_vector(15 downto 0);
    TILE0_RXUSRCLK0_IN                      : in   std_logic;
    TILE0_RXUSRCLK1_IN                      : in   std_logic;
    TILE0_RXUSRCLK20_IN                     : in   std_logic;
    TILE0_RXUSRCLK21_IN                     : in   std_logic;
    ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
    TILE0_RXN0_IN                           : in   std_logic;
    TILE0_RXN1_IN                           : in   std_logic;
    TILE0_RXP0_IN                           : in   std_logic;
    TILE0_RXP1_IN                           : in   std_logic;
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    TILE0_CLKIN_IN                          : in   std_logic;
    TILE0_GTPRESET_IN                       : in   std_logic;
    TILE0_PLLLKDET_OUT                      : out  std_logic;
    TILE0_REFCLKOUT_OUT                     : out  std_logic;
    TILE0_RESETDONE0_OUT                    : out  std_logic;
    TILE0_RESETDONE1_OUT                    : out  std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    TILE0_TXCHARISK0_IN                     : in   std_logic_vector(1 downto 0);
    TILE0_TXCHARISK1_IN                     : in   std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    TILE0_TXDATA0_IN                        : in   std_logic_vector(15 downto 0);
    TILE0_TXDATA1_IN                        : in   std_logic_vector(15 downto 0);
    TILE0_TXOUTCLK0_OUT                     : out  std_logic;
    TILE0_TXOUTCLK1_OUT                     : out  std_logic;
    TILE0_TXUSRCLK0_IN                      : in   std_logic;
    TILE0_TXUSRCLK1_IN                      : in   std_logic;
    TILE0_TXUSRCLK20_IN                     : in   std_logic;
    TILE0_TXUSRCLK21_IN                     : in   std_logic;
    --------------- Transmit Ports - TX Driver and OOB signalling --------------
    TILE0_TXN0_OUT                          : out  std_logic;
    TILE0_TXN1_OUT                          : out  std_logic;
    TILE0_TXP0_OUT                          : out  std_logic;
    TILE0_TXP1_OUT                          : out  std_logic


);
end component;


component MGT_USRCLK_SOURCE 
generic
(
    FREQUENCY_MODE   : string   := "LOW";    
    PERFORMANCE_MODE : string   := "MAX_SPEED"    
);
port
(
    DIV1_OUT                : out std_logic;
    DIV2_OUT                : out std_logic;
    DCM_LOCKED_OUT          : out std_logic;
    CLK_IN                  : in  std_logic;
    DCM_RESET_IN            : in  std_logic

);
end component;

component FRAME_GEN 
generic
(
    WORDS_IN_BRAM : integer    :=   256;
    MEM_00       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_01       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_02       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_03       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_04       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_05       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_06       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_07       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_08       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_09       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_10       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_11       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_12       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_13       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_14       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_15       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_16       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_17       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_18       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_19       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_20       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_21       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_22       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_23       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_24       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_25       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_26       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_27       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_28       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_29       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_30       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_31       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_32       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_33       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_34       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_35       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_36       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_37       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_38       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_39       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_00      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_01      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_02      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_03      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_04      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_05      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_06      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_07      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000"
);    
port
(
    -- User Interface
    TX_DATA             : out   std_logic_vector(31 downto 0);
    TX_CHARISK          : out   std_logic_vector(3 downto 0); 

    -- System Interface
    USER_CLK            : in    std_logic;
    SYSTEM_RESET        : in    std_logic
); 
end component;

component FRAME_CHECK 
generic
(
    RX_DATA_WIDTH            : integer := 16;
    USE_COMMA                : integer := 1;
    WORDS_IN_BRAM            : integer := 256;
    CONFIG_INDEPENDENT_LANES : integer := 0;
    START_OF_PACKET_CHAR     : std_logic_vector := x"55fb";
    MEM_00       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_01       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_02       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_03       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_04       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_05       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_06       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_07       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_08       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_09       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_0F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_10       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_11       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_12       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_13       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_14       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_15       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_16       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_17       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_18       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_19       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_1F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_20       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_21       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_22       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_23       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_24       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_25       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_26       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_27       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_28       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_29       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_2F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_30       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_31       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_32       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_33       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_34       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_35       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_36       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_37       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_38       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_39       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3A       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3B       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3C       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3D       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3E       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEM_3F       : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_00      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_01      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_02      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_03      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_04      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_05      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_06      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000";
    MEMP_07      : bit_vector :=   X"0000000000000000000000000000000000000000000000000000000000000000"
);
port
(
    -- User Interface
    RX_DATA                  : in  std_logic_vector((RX_DATA_WIDTH-1) downto 0); 
    RX_ENMCOMMA_ALIGN        : out std_logic;
    RX_ENPCOMMA_ALIGN        : out std_logic;
    RX_ENCHAN_SYNC           : out std_logic; 

    -- Control Interface
    INC_IN                   : in std_logic; 
    INC_OUT                  : out std_logic; 
    PATTERN_MATCH_N          : out std_logic;
    RESET_ON_ERROR           : in std_logic; 
    
    -- Error Monitoring
    ERROR_COUNT              : out std_logic_vector(7 downto 0);

    -- System Interface
    USER_CLK                 : in std_logic;
    SYSTEM_RESET             : in std_logic;
    TRACK_DATA               : out std_logic     
  
);
end component;

component MGT_USRCLK_SOURCE_PLL 
generic
(
    MULT                 : integer          := 2;
    DIVIDE               : integer          := 2;    
    CLK_PERIOD           : real             := 12.86;
    OUT0_DIVIDE          : integer          := 2;
    OUT1_DIVIDE          : integer          := 2;
    OUT2_DIVIDE          : integer          := 2;
    OUT3_DIVIDE          : integer          := 2;
    SIMULATION_P         : integer          := 1;
    LOCK_WAIT_COUNT      : std_logic_vector := "1000001000110101"    
);
port
( 
    CLK0_OUT                : out std_logic;
    CLK1_OUT                : out std_logic;
    CLK2_OUT                : out std_logic;
    CLK3_OUT                : out std_logic;
    CLK_IN                  : in  std_logic;
    PLL_LOCKED_OUT          : out std_logic;
    PLL_RESET_IN            : in  std_logic
);
end component;





-- Chipscope modules
attribute syn_black_box                : boolean;
attribute syn_noprune                  : boolean;


component shared_vio
port
(
    control                 : in  std_logic_vector(35 downto 0);
    async_in                : in  std_logic_vector(31 downto 0);
    async_out               : out std_logic_vector(31 downto 0)
);
end component;
attribute syn_black_box of shared_vio : component is TRUE;
attribute syn_noprune of shared_vio   : component is TRUE;


component icon
port
(
    control0                : out std_logic_vector(35 downto 0);
    control1                : out std_logic_vector(35 downto 0);
    control2                : out std_logic_vector(35 downto 0);
    control3                : out std_logic_vector(35 downto 0);
    control4                : out std_logic_vector(35 downto 0);
    control5                : out std_logic_vector(35 downto 0);
    control6                : out std_logic_vector(35 downto 0)
);
end component;
attribute syn_black_box of icon : component is TRUE;
attribute syn_noprune of icon   : component is TRUE;


component ila
port
(
    control                 : in  std_logic_vector(35 downto 0);
    clk                     : in  std_logic;
    trig0                   : in  std_logic_vector(63 downto 0)
);
end component;
attribute syn_black_box of ila : component is TRUE;
attribute syn_noprune of ila   : component is TRUE;


--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;
    
--************************** Register Declarations ****************************

    signal     tile0_tx_resetdone0_r           : std_logic;
    signal     tile0_tx_resetdone0_r2          : std_logic;
    signal     tile0_tx_resetdone1_r           : std_logic;
    signal     tile0_tx_resetdone1_r2          : std_logic;
    signal     tile0_rx_resetdone0_r           : std_logic;
    signal     tile0_rx_resetdone0_r2          : std_logic;
    signal     tile0_rx_resetdone1_r           : std_logic;
    signal     tile0_rx_resetdone1_r2          : std_logic;
 
    

--**************************** Wire Declarations ******************************

    -------------------------- MGT Wrapper Wires ------------------------------
    --________________________________________________________________________
    --________________________________________________________________________
    --TILE0   (X0Y5)

    ----------------------- Receive Ports - 8b10b Decoder ----------------------
    signal  tile0_rxchariscomma0_i          : std_logic_vector(1 downto 0);
    signal  tile0_rxchariscomma1_i          : std_logic_vector(1 downto 0);
    signal  tile0_rxcharisk0_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxcharisk1_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxdisperr0_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxdisperr1_i              : std_logic_vector(1 downto 0);
    signal  tile0_rxnotintable0_i           : std_logic_vector(1 downto 0);
    signal  tile0_rxnotintable1_i           : std_logic_vector(1 downto 0);
    --------------- Receive Ports - Comma Detection and Alignment --------------
    signal  tile0_rxbyteisaligned0_i        : std_logic;
    signal  tile0_rxbyteisaligned1_i        : std_logic;
    signal  tile0_rxenmcommaalign0_i        : std_logic;
    signal  tile0_rxenmcommaalign1_i        : std_logic;
    signal  tile0_rxenpcommaalign0_i        : std_logic;
    signal  tile0_rxenpcommaalign1_i        : std_logic;
    ------------------- Receive Ports - RX Data Path interface -----------------
    signal  tile0_rxdata0_i                 : std_logic_vector(15 downto 0);
    signal  tile0_rxdata1_i                 : std_logic_vector(15 downto 0);
    --------------------- Shared Ports - Tile and PLL Ports --------------------
    signal  tile0_gtpreset_i                : std_logic;
    signal  tile0_plllkdet_i                : std_logic;
    signal  tile0_refclkout_i               : std_logic;
    signal  tile0_resetdone0_i              : std_logic;
    signal  tile0_resetdone1_i              : std_logic;
    ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
    signal  tile0_txcharisk0_i              : std_logic_vector(1 downto 0);
    signal  tile0_txcharisk1_i              : std_logic_vector(1 downto 0);
    ------------------ Transmit Ports - TX Data Path interface -----------------
    signal  tile0_txdata0_i                 : std_logic_vector(15 downto 0);
    signal  tile0_txdata1_i                 : std_logic_vector(15 downto 0);
    signal  tile0_txoutclk0_i               : std_logic;
    signal  tile0_txoutclk1_i               : std_logic;


    ------------------------------- Global Signals -----------------------------
    signal  tile0_tx_system_reset0_c        : std_logic;
    signal  tile0_rx_system_reset0_c        : std_logic;
    signal  tile0_rxreset0_i                : std_logic;
    signal  tile0_txreset0_i                : std_logic;
    signal  tile0_tx_system_reset1_c        : std_logic;
    signal  tile0_rx_system_reset1_c        : std_logic;
    signal  tile0_rxreset1_i                : std_logic;
    signal  tile0_txreset1_i                : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drp_clk_in_i                    : std_logic;
    signal  tile0_refclkout_bufg_i          : std_logic;
    
    
    ----------------------------- User Clocks ---------------------------------
    signal  tile0_txusrclk0_i               : std_logic;
    signal  tile0_txusrclk20_i              : std_logic;
    signal  refclkout_pll0_locked_i         : std_logic;
    signal  refclkout_pll0_reset_i          : std_logic;
    signal  tile0_refclkout_to_cmt_i        : std_logic;


    ----------------------- Frame check/gen Module Signals --------------------
    signal  tile0_refclk_i                  : std_logic;
    signal  tile0_matchn0_i                 : std_logic;
    signal  tile0_track_data0_i             : std_logic;    
    signal  tile0_txcharisk0_float_i        : std_logic_vector(1 downto 0);
    signal  tile0_txdata0_float_i           : std_logic_vector(15 downto 0);
    signal  tile0_error_count0_i            : std_logic_vector(7 downto 0);
    signal  tile0_frame_check0_reset_i      : std_logic;
    signal  tile0_inc_in0_i                 : std_logic;
    signal  tile0_inc_out0_i                : std_logic;
    signal  tile0_matchn1_i                 : std_logic;
    signal  tile0_track_data1_i             : std_logic;    
    signal  tile0_txcharisk1_float_i        : std_logic_vector(1 downto 0);
    signal  tile0_txdata1_float_i           : std_logic_vector(15 downto 0);
    signal  tile0_error_count1_i            : std_logic_vector(7 downto 0);
    signal  tile0_frame_check1_reset_i      : std_logic;
    signal  tile0_inc_in1_i                 : std_logic;
    signal  tile0_inc_out1_i                : std_logic;

    signal  reset_on_data_error_i           : std_logic;
    
    ------------------------- Sync Module Signals -----------------------------
    signal  tx_sync_done_i                  : std_logic;
    
    signal  reset_txsync_c                  : std_logic;
    signal    track_data_out_i                : std_logic;

    ----------------------- Chipscope Signals ---------------------------------

    signal  shared_vio_control_i            : std_logic_vector(35 downto 0);
    signal  tx_data_vio_control0_i          : std_logic_vector(35 downto 0);
    signal  rx_data_vio_control0_i          : std_logic_vector(35 downto 0);
    signal  ila_control0_i                  : std_logic_vector(35 downto 0);
    signal  tx_data_vio_control1_i          : std_logic_vector(35 downto 0);
    signal  rx_data_vio_control1_i          : std_logic_vector(35 downto 0);
    signal  ila_control1_i                  : std_logic_vector(35 downto 0);
    signal  shared_vio_in_i                 : std_logic_vector(31 downto 0);
    signal  shared_vio_out_i                : std_logic_vector(31 downto 0);
    signal  tx_data_vio_in0_i               : std_logic_vector(31 downto 0);
    signal  tx_data_vio_out0_i              : std_logic_vector(31 downto 0);
    signal  tx_data_vio_in1_i               : std_logic_vector(31 downto 0);
    signal  tx_data_vio_out1_i              : std_logic_vector(31 downto 0);
    signal  rx_data_vio_in0_i               : std_logic_vector(31 downto 0);
    signal  rx_data_vio_out0_i              : std_logic_vector(31 downto 0);
    signal  rx_data_vio_in1_i               : std_logic_vector(31 downto 0);
    signal  rx_data_vio_out1_i              : std_logic_vector(31 downto 0);
    signal  ila_in0_i                       : std_logic_vector(63 downto 0);
    signal  ila_in1_i                       : std_logic_vector(63 downto 0);

    signal  tile0_tx_data_vio_in0_i         : std_logic_vector(31 downto 0);
    signal  tile0_tx_data_vio_out0_i        : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_in0_i         : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_out0_i        : std_logic_vector(31 downto 0);
    signal  tile0_ila_in0_i                 : std_logic_vector(63 downto 0);
    signal  tile0_tx_data_vio_in1_i         : std_logic_vector(31 downto 0);
    signal  tile0_tx_data_vio_out1_i        : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_in1_i         : std_logic_vector(31 downto 0);
    signal  tile0_rx_data_vio_out1_i        : std_logic_vector(31 downto 0);
    signal  tile0_ila_in1_i                 : std_logic_vector(63 downto 0);


    signal  gtpreset_i                      : std_logic;
    signal  user_tx_reset_i                 : std_logic;
    signal  user_rx_reset_i                 : std_logic;
    signal  ila_clk0_i                      : std_logic;
    signal  ila_clk_mux_out0_i              : std_logic;
    signal  ila_clk1_i                      : std_logic;
    signal  ila_clk_mux_out1_i              : std_logic;


--**************************** Main Body of Code *******************************
begin

    --  Static signal Assigments
    tied_to_ground_i                        <= '0';
    tied_to_ground_vec_i                    <= x"0000000000000000";
    tied_to_vcc_i                           <= '1';
    tied_to_vcc_vec_i                       <= x"ff";


    


    -----------------------Dedicated GTP Reference Clock Inputs ---------------
    -- The dedicated reference clock inputs you selected in the GUI are implemented using
    -- IBUFDS instances.
    --
    -- In the UCF file for this example design, you will see that each of
    -- these IBUFDS instances has been LOCed to a particular set of pins. By LOCing to these
    -- locations, we tell the tools to use the dedicated input buffers to the GTP reference
    -- clock network, rather than general purpose IOs. To select other pins, consult the 
    -- Implementation chapter of UG196, or rerun the wizard.
    --
    -- This network is the highest performace (lowest jitter) option for providing clocks
    -- to the GTP transceivers.
    
    tile0_refclk_ibufds_i : IBUFDS
    port map
    (
        O                               =>      tile0_refclk_i,
        I                               =>      TILE0_REFCLK_PAD_P_IN,
        IB                              =>      TILE0_REFCLK_PAD_N_IN
    );






    ----------------------------------- User Clocks ---------------------------
    
    -- The clock resources in this section were added based on userclk source selections on
    -- the Latency, Buffering, and Clocking page of the GUI. A few notes about user clocks:
    -- * The userclk and userclk2 for each GTP datapath (TX and RX) must be phase aligned to 
    --   avoid data errors in the fabric interface whenever the datapath is wider than 10 bits
    -- * To minimize clock resources, you can share clocks between GTPs. GTPs using the same frequency
    --   or multiples of the same frequency can be accomadated using DCMs and PLLs. Use caution when
    --   using RXRECCLK as a clock source, however - these clocks can typically only be shared if all
    --   the channels using the clock are receiving data from TX channels that share a reference clock 
    --   source with each other.

    refclkout_pll0_bufg_i : BUFG
    port map
    (
        I                               =>      tile0_refclkout_i,
        O                               =>      tile0_refclkout_to_cmt_i
    );

    refclkout_pll0_reset_i                  <= not tile0_plllkdet_i;
    refclkout_pll0_i : MGT_USRCLK_SOURCE_PLL
    generic map
    (
        MULT                            =>      10,
        DIVIDE                          =>      1,
        CLK_PERIOD                      =>      12.86,
        OUT0_DIVIDE                     =>      10,
        OUT1_DIVIDE                     =>      5,
        OUT2_DIVIDE                     =>      1,
        OUT3_DIVIDE                     =>      1,
        SIMULATION_P                    =>      EXAMPLE_USE_CHIPSCOPE,
        LOCK_WAIT_COUNT                 =>      "0001111001100000"
    )
    port map
    (
        CLK0_OUT                        =>      tile0_txusrclk20_i,
        CLK1_OUT                        =>      tile0_txusrclk0_i,
        CLK2_OUT                        =>      open,
        CLK3_OUT                        =>      open,
        CLK_IN                          =>      tile0_refclkout_to_cmt_i,
        PLL_LOCKED_OUT                  =>      refclkout_pll0_locked_i,
        PLL_RESET_IN                    =>      refclkout_pll0_reset_i
    );






    ----------------------------- The GTP Wrapper -----------------------------
    
    -- Use the instantiation template in the project directory to add the GTP wrapper to your design.
    -- In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    -- checker. The GTPs will reset, then attempt to align and transmit data. If channel bonding is 
    -- enabled, bonding should occur after alignment.
    

    -- Wire all PLLLKDET signals to the top level as output ports
    TILE0_PLLLKDET_OUT                      <= tile0_plllkdet_i;



    single_channel_aurora_xc5vsx95t_i : SINGLE_CHANNEL_AURORA_XC5VSX95T
    generic map
    (
        WRAPPER_SIM_MODE                =>      EXAMPLE_SIM_MODE,   
        WRAPPER_SIM_GTPRESET_SPEEDUP    =>      EXAMPLE_SIM_GTPRESET_SPEEDUP,
        WRAPPER_SIM_PLL_PERDIV2         =>      EXAMPLE_SIM_PLL_PERDIV2
    )
    port map
    (
    
 
 
 
 

 
 
 
 

        --_____________________________________________________________________
        --_____________________________________________________________________
        --TILE0  (X0Y5)

        ----------------------- Receive Ports - 8b10b Decoder ----------------------
        TILE0_RXCHARISCOMMA0_OUT        =>      tile0_rxchariscomma0_i,
        TILE0_RXCHARISCOMMA1_OUT        =>      tile0_rxchariscomma1_i,
        TILE0_RXCHARISK0_OUT            =>      tile0_rxcharisk0_i,
        TILE0_RXCHARISK1_OUT            =>      tile0_rxcharisk1_i,
        TILE0_RXDISPERR0_OUT            =>      tile0_rxdisperr0_i,
        TILE0_RXDISPERR1_OUT            =>      tile0_rxdisperr1_i,
        TILE0_RXNOTINTABLE0_OUT         =>      tile0_rxnotintable0_i,
        TILE0_RXNOTINTABLE1_OUT         =>      tile0_rxnotintable1_i,
        --------------- Receive Ports - Comma Detection and Alignment --------------
        TILE0_RXBYTEISALIGNED0_OUT      =>      tile0_rxbyteisaligned0_i,
        TILE0_RXBYTEISALIGNED1_OUT      =>      tile0_rxbyteisaligned1_i,
        TILE0_RXENMCOMMAALIGN0_IN       =>      tile0_rxenmcommaalign0_i,
        TILE0_RXENMCOMMAALIGN1_IN       =>      tile0_rxenmcommaalign1_i,
        TILE0_RXENPCOMMAALIGN0_IN       =>      tile0_rxenpcommaalign0_i,
        TILE0_RXENPCOMMAALIGN1_IN       =>      tile0_rxenpcommaalign1_i,
        ------------------- Receive Ports - RX Data Path interface -----------------
        TILE0_RXDATA0_OUT               =>      tile0_rxdata0_i,
        TILE0_RXDATA1_OUT               =>      tile0_rxdata1_i,
        TILE0_RXUSRCLK0_IN              =>      tile0_txusrclk0_i,
        TILE0_RXUSRCLK1_IN              =>      tile0_txusrclk0_i,
        TILE0_RXUSRCLK20_IN             =>      tile0_txusrclk20_i,
        TILE0_RXUSRCLK21_IN             =>      tile0_txusrclk20_i,
        ------- Receive Ports - RX Driver,OOB signalling,Coupling and Eq.,CDR ------
        TILE0_RXN0_IN                   =>      RXN_IN(0),
        TILE0_RXN1_IN                   =>      RXN_IN(1),
        TILE0_RXP0_IN                   =>      RXP_IN(0),
        TILE0_RXP1_IN                   =>      RXP_IN(1),
        --------------------- Shared Ports - Tile and PLL Ports --------------------
        TILE0_CLKIN_IN                  =>      tile0_refclk_i,
        TILE0_GTPRESET_IN               =>      tile0_gtpreset_i,
        TILE0_PLLLKDET_OUT              =>      tile0_plllkdet_i,
        TILE0_REFCLKOUT_OUT             =>      tile0_refclkout_i,
        TILE0_RESETDONE0_OUT            =>      tile0_resetdone0_i,
        TILE0_RESETDONE1_OUT            =>      tile0_resetdone1_i,
        ---------------- Transmit Ports - 8b10b Encoder Control Ports --------------
        TILE0_TXCHARISK0_IN             =>      tile0_txcharisk0_i,
        TILE0_TXCHARISK1_IN             =>      tile0_txcharisk1_i,
        ------------------ Transmit Ports - TX Data Path interface -----------------
        TILE0_TXDATA0_IN                =>      tile0_txdata0_i,
        TILE0_TXDATA1_IN                =>      tile0_txdata1_i,
        TILE0_TXOUTCLK0_OUT             =>      tile0_txoutclk0_i,
        TILE0_TXOUTCLK1_OUT             =>      tile0_txoutclk1_i,
        TILE0_TXUSRCLK0_IN              =>      tile0_txusrclk0_i,
        TILE0_TXUSRCLK1_IN              =>      tile0_txusrclk0_i,
        TILE0_TXUSRCLK20_IN             =>      tile0_txusrclk20_i,
        TILE0_TXUSRCLK21_IN             =>      tile0_txusrclk20_i,
        --------------- Transmit Ports - TX Driver and OOB signalling --------------
        TILE0_TXN0_OUT                  =>      TXN_OUT(0),
        TILE0_TXN1_OUT                  =>      TXN_OUT(1),
        TILE0_TXP0_OUT                  =>      TXP_OUT(0),
        TILE0_TXP1_OUT                  =>      TXP_OUT(1)


    );






    -------------------------- User Module Resets -----------------------------
    -- All the User Modules i.e. FRAME_GEN, FRAME_CHECK and the sync modules
    -- are held in reset till the RESETDONE goes high. 
    -- The RESETDONE is registered a couple of times on USRCLK2 and connected 
    -- to the reset of the modules
    
    process( tile0_txusrclk20_i,tile0_resetdone0_i)
    begin
        if(tile0_resetdone0_i = '0') then
            tile0_rx_resetdone0_r  <= '0'   after DLY;
            tile0_rx_resetdone0_r2 <= '0'   after DLY;
        elsif(tile0_txusrclk20_i'event and tile0_txusrclk20_i = '1') then
            tile0_rx_resetdone0_r  <= tile0_resetdone0_i   after DLY;
            tile0_rx_resetdone0_r2 <= tile0_rx_resetdone0_r   after DLY;
        end if;
    end process;
    
    process( tile0_txusrclk20_i,tile0_resetdone1_i)
    begin
        if(tile0_resetdone1_i = '0') then
            tile0_rx_resetdone1_r  <= '0'   after DLY;
            tile0_rx_resetdone1_r2 <= '0'   after DLY;
        elsif(tile0_txusrclk20_i'event and tile0_txusrclk20_i = '1') then
            tile0_rx_resetdone1_r  <= tile0_resetdone1_i   after DLY;
            tile0_rx_resetdone1_r2 <= tile0_rx_resetdone1_r   after DLY;
        end if;
    end process;
    
    process( tile0_txusrclk20_i,tile0_resetdone0_i)
    begin
        if (tile0_resetdone0_i = '0') then 
            tile0_tx_resetdone0_r    <=   '0'	after DLY ;
            tile0_tx_resetdone0_r2   <=   '0'	after DLY ;
        elsif(tile0_txusrclk20_i'event and tile0_txusrclk20_i = '1') then
            tile0_tx_resetdone0_r    <=   tile0_resetdone0_i	after DLY;
            tile0_tx_resetdone0_r2   <=   tile0_tx_resetdone0_r	after DLY;
        end if;
    end process; 
    process( tile0_txusrclk20_i,tile0_resetdone1_i)
    begin
        if (tile0_resetdone1_i = '0') then 
            tile0_tx_resetdone1_r    <=   '0'	after DLY ;
            tile0_tx_resetdone1_r2   <=   '0'	after DLY ;
        elsif(tile0_txusrclk20_i'event and tile0_txusrclk20_i = '1') then
            tile0_tx_resetdone1_r    <=   tile0_resetdone1_i	after DLY;
            tile0_tx_resetdone1_r2   <=   tile0_tx_resetdone1_r	after DLY;
        end if;
    end process; 
    



    ------------------------------ Frame Generators ---------------------------
    -- The example design uses Block RAM based frame generators to provide test
    -- data to the GTPs for transmission. By default the frame generators are 
    -- loaded with an incrementing data sequence that includes commas/alignment
    -- characters for alignment. If your protocol uses channel bonding, the 
    -- frame generator will also be preloaded with a channel bonding sequence.
    
    -- You can modify the data transmitted by changing the INIT values of the frame
    -- generator in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.

    tile0_frame_gen0 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_01                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_02                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_03                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_04                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_05                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_06                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_07                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_08                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_09                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_0A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_0B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_0C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_0D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_0E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_0F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_10                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_11                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_12                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_13                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_14                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_15                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_16                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_17                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_18                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_19                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_1A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_1B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_1C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_1D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_1E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_1F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_20                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_21                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_22                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_23                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_24                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_25                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_26                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_27                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_28                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_29                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_2A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_2B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_2C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_2D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_2E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_2F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_30                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_31                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_32                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_33                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_34                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_35                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_36                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_37                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_38                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_39                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_3A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_3B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_3C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_3D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_3E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_3F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000003"
    )
    port map
    (
        -- User Interface
        TX_DATA(31 downto 16)           =>      tile0_txdata0_float_i,
        TX_DATA(15 downto 0)            =>      tile0_txdata0_i,
        TX_CHARISK(3 downto 2)          =>      tile0_txcharisk0_float_i,
        TX_CHARISK(1 downto 0)          =>      tile0_txcharisk0_i,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk20_i,
        SYSTEM_RESET                    =>      tile0_tx_system_reset0_c
    );
    
    tile0_frame_gen1 : FRAME_GEN
    generic map
    (
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        MEM_00                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_01                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_02                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_03                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_04                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_05                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_06                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_07                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_08                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_09                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_0A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_0B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_0C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_0D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_0E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_0F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_10                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_11                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_12                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_13                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_14                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_15                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_16                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_17                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_18                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_19                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_1A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_1B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_1C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_1D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_1E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_1F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_20                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_21                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_22                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_23                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_24                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_25                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_26                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_27                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_28                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_29                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_2A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_2B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_2C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_2D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_2E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_2F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_30                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_31                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_32                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_33                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_34                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_35                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_36                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_37                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_38                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_39                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_3A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_3B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_3C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_3D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_3E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_3F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000003"
    )
    port map
    (
        -- User Interface
        TX_DATA(31 downto 16)           =>      tile0_txdata1_float_i,
        TX_DATA(15 downto 0)            =>      tile0_txdata1_i,
        TX_CHARISK(3 downto 2)          =>      tile0_txcharisk1_float_i,
        TX_CHARISK(1 downto 0)          =>      tile0_txcharisk1_i,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk20_i,
        SYSTEM_RESET                    =>      tile0_tx_system_reset1_c
    );
    


    ---------------------------------- Frame Checkers -------------------------
    -- The example design uses Block RAM based frame checkers to verify incoming  
    -- data. By default the frame generators are loaded with a data sequence that 
    -- matches the outgoing sequence of the frame generators for the TX ports.
    
    -- You can modify the expected data sequence by changing the INIT values of the frame
    -- checkers in this file. Pay careful attention to bit order and the spacing
    -- of your control and alignment characters.
    
    -- When the frame checker receives data, it attempts to synchronise to the 
    -- incoming pattern by looking for the first sequence in the pattern. Once it 
    -- finds the first sequence, it increments through the sequence, and indicates an 
    -- error whenever the next value received does not match the expected value.

    tile0_frame_check0_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile0_matchn0_i;

    -- tile0_frame_check0 is always connected to the lane with the start of char
    -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    tile0_inc_in0_i                         <= '0';

    tile0_frame_check0 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      1,
        START_OF_PACKET_CHAR            =>      x"bcbc",
        MEM_00                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_01                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_02                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_03                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_04                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_05                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_06                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_07                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_08                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_09                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_0A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_0B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_0C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_0D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_0E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_0F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_10                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_11                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_12                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_13                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_14                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_15                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_16                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_17                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_18                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_19                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_1A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_1B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_1C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_1D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_1E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_1F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_20                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_21                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_22                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_23                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_24                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_25                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_26                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_27                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_28                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_29                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_2A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_2B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_2C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_2D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_2E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_2F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_30                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_31                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_32                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_33                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_34                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_35                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_36                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_37                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_38                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_39                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_3A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_3B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_3C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_3D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_3E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_3F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000003"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile0_rxdata0_i,
        RX_ENMCOMMA_ALIGN               =>      tile0_rxenmcommaalign0_i,
        RX_ENPCOMMA_ALIGN               =>      tile0_rxenpcommaalign0_i,
        RX_ENCHAN_SYNC                  =>      open,
        -- Control Interface
        INC_IN                          =>      tile0_inc_in0_i,
        INC_OUT                         =>      tile0_inc_out0_i,
        PATTERN_MATCH_N                 =>      tile0_matchn0_i,
        RESET_ON_ERROR                  =>      tile0_frame_check0_reset_i,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk20_i,
        SYSTEM_RESET                    =>      tile0_rx_system_reset0_c,
        ERROR_COUNT                     =>      tile0_error_count0_i,
        TRACK_DATA                      =>      tile0_track_data0_i
    );
    
    tile0_frame_check1_reset_i              <= reset_on_data_error_i when (EXAMPLE_CONFIG_INDEPENDENT_LANES=0) else tile0_matchn1_i;

    -- tile0_frame_check0 is always connected to the lane with the start of char
    -- and this lane starts off the data checking on all the other lanes. The INC_IN port is tied off
    tile0_inc_in1_i                         <= '0';

    tile0_frame_check1 : FRAME_CHECK
    generic map
    (
        RX_DATA_WIDTH                   =>      16,
        USE_COMMA                       =>      1,
        WORDS_IN_BRAM                   =>      EXAMPLE_WORDS_IN_BRAM,
        CONFIG_INDEPENDENT_LANES        =>      1,
        START_OF_PACKET_CHAR            =>      x"bcbc",
        MEM_00                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_01                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_02                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_03                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_04                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_05                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_06                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_07                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_08                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_09                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_0A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_0B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_0C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_0D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_0E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_0F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_10                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_11                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_12                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_13                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_14                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_15                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_16                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_17                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_18                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_19                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_1A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_1B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_1C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_1D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_1E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_1F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_20                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_21                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_22                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_23                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_24                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_25                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_26                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_27                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_28                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_29                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_2A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_2B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_2C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_2D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_2E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_2F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_30                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_31                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_32                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_33                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_34                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_35                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_36                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_37                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEM_38                  =>  x"00000d0c00000b0a00000908000007060000050400000302000001000000bcbc",
        MEM_39                  =>  x"00001d1c00001b1a000019180000171600001514000013120000111000000f0e",
        MEM_3A                  =>  x"00002d2c00002b2a000029280000272600002524000023220000212000001f1e",
        MEM_3B                  =>  x"00003d3c00003b3a000039380000373600003534000033320000313000002f2e",
        MEM_3C                  =>  x"00004d4c00004b4a000049480000474600004544000043420000414000003f3e",
        MEM_3D                  =>  x"00005d5c00005b5a000059580000575600005554000053520000515000004f4e",
        MEM_3E                  =>  x"00006d6c00006b6a000069680000676600006564000063620000616000005f5e",
        MEM_3F                  =>  x"00007d7c00007b7a000079780000777600007574000073720000717000006f6e",
        MEMP_00                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_01                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_02                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_03                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_04                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_05                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_06                  =>  x"0000000000000000000000000000000000000000000000000000000000000003",
        MEMP_07                  =>  x"0000000000000000000000000000000000000000000000000000000000000003"
    )
    port map
    (
        -- MGT Interface
        RX_DATA                         =>      tile0_rxdata1_i,
        RX_ENMCOMMA_ALIGN               =>      tile0_rxenmcommaalign1_i,
        RX_ENPCOMMA_ALIGN               =>      tile0_rxenpcommaalign1_i,
        RX_ENCHAN_SYNC                  =>      open,
        -- Control Interface
        INC_IN                          =>      tile0_inc_in1_i,
        INC_OUT                         =>      tile0_inc_out1_i,
        PATTERN_MATCH_N                 =>      tile0_matchn1_i,
        RESET_ON_ERROR                  =>      tile0_frame_check1_reset_i,
        -- System Interface
        USER_CLK                        =>      tile0_txusrclk20_i,
        SYSTEM_RESET                    =>      tile0_rx_system_reset1_c,
        ERROR_COUNT                     =>      tile0_error_count1_i,
        TRACK_DATA                      =>      tile0_track_data1_i
    );
    



    TRACK_DATA_OUT                          <= track_data_out_i;
    
    track_data_out_i                        <= 
                                tile0_track_data0_i and
                                tile0_track_data1_i 
 ;

    ----------------------------- Chipscope Connections -----------------------
    -- When the example design is run in hardware, it uses chipscope to allow the
    -- example design and GTP wrapper to be controlled and monitored. The 
    -- EXAMPLE_USE_CHIPSCOPE parameter allows chipscope to be removed for simulation.
    
chipscope : if EXAMPLE_USE_CHIPSCOPE = 1 generate


    -- Shared VIO for all tiles
    shared_vio_i : shared_vio
    port map
    (
        control                         =>      shared_vio_control_i,
        async_in                        =>      shared_vio_in_i,
        async_out                       =>      shared_vio_out_i
    );

    
    -- ICON for all VIOs 
    i_icon : icon
    port map
    (
        control0                        =>      shared_vio_control_i,
        control1                        =>      tx_data_vio_control0_i,
        control2                        =>      rx_data_vio_control0_i,
        control3                        =>      ila_control0_i,
        control4                        =>      tx_data_vio_control1_i,
        control5                        =>      rx_data_vio_control1_i,
        control6                        =>      ila_control1_i
    );

    -- TX VIO 
    tx_data_vio0_i : shared_vio
    port map
    (
        control                         =>      tx_data_vio_control0_i,
        async_in                        =>      tx_data_vio_in0_i,
        async_out                       =>      tx_data_vio_out0_i
    );
    
    -- RX VIO 
    rx_data_vio0_i : shared_vio
    port map
    (
        control                         =>      rx_data_vio_control0_i,
        async_in                        =>      rx_data_vio_in0_i,
        async_out                       =>      rx_data_vio_out0_i
    );
    
    -- RX ILA
    ila0_i : ila
    port map
    (
        control                         =>      ila_control0_i,
        clk                             =>      ila_clk0_i,
        trig0                           =>      ila_in0_i
    );

    -- The RX ILA must use the same clock as the selected transceiver
    ila_clk0_bufg_i : BUFG
    port map
    (
        I => ila_clk_mux_out0_i,
        O => ila_clk0_i
    );

     ila_clk_mux_out0_i<= tile0_txusrclk20_i;

        
    -- TX VIO 
    tx_data_vio1_i : shared_vio
    port map
    (
        control                         =>      tx_data_vio_control1_i,
        async_in                        =>      tx_data_vio_in1_i,
        async_out                       =>      tx_data_vio_out1_i
    );
    
    -- RX VIO 
    rx_data_vio1_i : shared_vio
    port map
    (
        control                         =>      rx_data_vio_control1_i,
        async_in                        =>      rx_data_vio_in1_i,
        async_out                       =>      rx_data_vio_out1_i
    );
    
    -- RX ILA
    ila1_i : ila
    port map
    (
        control                         =>      ila_control1_i,
        clk                             =>      ila_clk1_i,
        trig0                           =>      ila_in1_i
    );

    -- The RX ILA must use the same clock as the selected transceiver
    ila_clk1_bufg_i : BUFG
    port map
    (
        I => ila_clk_mux_out1_i,
        O => ila_clk1_i
    );

     ila_clk_mux_out1_i<= tile0_txusrclk20_i;

        

    -- Connect resets for frame generators
    tile0_tx_system_reset0_c                <= not tile0_tx_resetdone0_r2 or user_tx_reset_i;
    tile0_tx_system_reset1_c                <= not tile0_tx_resetdone1_r2 or user_tx_reset_i;
    tile0_rx_system_reset0_c                <= not tile0_rx_resetdone0_r2 or user_rx_reset_i;
    tile0_rx_system_reset1_c                <= not tile0_rx_resetdone1_r2 or user_rx_reset_i;


    tile0_gtpreset_i                        <= gtpreset_i;


    -- Shared VIO Outputs
    gtpreset_i                              <= shared_vio_out_i(31);
    user_tx_reset_i                         <= shared_vio_out_i(30);
    user_rx_reset_i                         <= shared_vio_out_i(29);

    -- Shared VIO Inputs
    shared_vio_in_i(31)                     <= tile0_plllkdet_i;
    shared_vio_in_i(30 downto 0)            <= "0000000000000000000000000000000";

    -- Chipscope connections for GTP0 on Tile 0
    tile0_tx_data_vio_in0_i(31 downto 0)    <= "00000000000000000000000000000000";
    tile0_rx_data_vio_in0_i(31)             <= tile0_resetdone0_i;
    tile0_rx_data_vio_in0_i(30 downto 0)    <= "0000000000000000000000000000000";
    tile0_ila_in0_i(63 downto 62)           <= tile0_rxchariscomma0_i;
    tile0_ila_in0_i(61 downto 60)           <= tile0_rxcharisk0_i;
    tile0_ila_in0_i(59 downto 58)           <= tile0_rxdisperr0_i;
    tile0_ila_in0_i(57 downto 56)           <= tile0_rxnotintable0_i;
    tile0_ila_in0_i(55)                     <= tile0_rxbyteisaligned0_i;
    tile0_ila_in0_i(54 downto 39)           <= tile0_rxdata0_i;
    tile0_ila_in0_i(38 downto 31)           <= tile0_error_count0_i;
    tile0_ila_in0_i(30 downto 0)            <= "0000000000000000000000000000000";

    -- Chipscope connections for GTP1 on Tile 0
    tile0_tx_data_vio_in1_i(31 downto 0)    <= "00000000000000000000000000000000";
    tile0_rx_data_vio_in1_i(31)             <= tile0_resetdone1_i;
    tile0_rx_data_vio_in1_i(30 downto 0)    <= "0000000000000000000000000000000";
    tile0_ila_in1_i(63 downto 62)           <= tile0_rxchariscomma1_i;
    tile0_ila_in1_i(61 downto 60)           <= tile0_rxcharisk1_i;
    tile0_ila_in1_i(59 downto 58)           <= tile0_rxdisperr1_i;
    tile0_ila_in1_i(57 downto 56)           <= tile0_rxnotintable1_i;
    tile0_ila_in1_i(55)                     <= tile0_rxbyteisaligned1_i;
    tile0_ila_in1_i(54 downto 39)           <= tile0_rxdata1_i;
    tile0_ila_in1_i(38 downto 31)           <= tile0_error_count1_i;
    tile0_ila_in1_i(30 downto 0)            <= "0000000000000000000000000000000";


    tx_data_vio_in0_i                   <=      tile0_tx_data_vio_in0_i;


    rx_data_vio_in0_i                   <=      tile0_rx_data_vio_in0_i;


    ila_in0_i                           <=      tile0_ila_in0_i;


    tx_data_vio_in1_i                   <=      tile0_tx_data_vio_in1_i;


    rx_data_vio_in1_i                   <=      tile0_rx_data_vio_in1_i;


    ila_in1_i                           <=      tile0_ila_in1_i;




   
end generate chipscope;


no_chipscope : if EXAMPLE_USE_CHIPSCOPE = 0 generate

    -- If Chipscope is not being used, drive GTP reset signal
    -- from the top level ports
    tile0_gtpreset_i                        <= GTPRESET_IN;

    -- assign resets for frame_gen and frame_check modules
    tile0_tx_system_reset0_c                <= not tile0_tx_resetdone0_r2;
    tile0_tx_system_reset1_c                <= not tile0_tx_resetdone1_r2;
    tile0_rx_system_reset0_c                <= not tile0_rx_resetdone0_r2;
    tile0_rx_system_reset1_c                <= not tile0_rx_resetdone1_r2;



    gtpreset_i                              <= tied_to_ground_i;
    user_tx_reset_i                         <= tied_to_ground_i;
    user_rx_reset_i                         <= tied_to_ground_i;



end generate no_chipscope;


end RTL;

